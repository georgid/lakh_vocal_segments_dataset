BZh91AY&SYt�aa_�ryg����������`�^� �;wYA�����eS��:�`ٶѭi���[7]�@۶�q�;��n\wx |E ET@  $U  M�E�lR��4
�T4"�����( �Ǩ!��B�/��:�+��:n�l0����{t�XH[8��Q��z m��n��
��6�w���'�U.��C��Z�C�i�]��@	[�т��|�L��^�;�tzu�F�`!�Z�]�����n�)v���h��-����M�;9Ev���((/�*�i�w`�m�[��!��I��O�F�:�xt�`PPm�JࠣϽ�q�(o:�pS�A���T�dC��|X��T�R���PPm�}�9:4BeQ����w$��׻�ފW��;�PHm�Ҹ(���(;��ǔ�  }Q����W�A�|��.
0Pd��(n�*࠶p�
��彆 AA��4�+�[}�9)"�R�
�P�(�TU
�!��#OT�J���&� �# & ����=U*�@         ��UJ552����@C  ���T���P�4h  ��  *	@�4%?M5O�M�OT?H�z�S�z��4�
�)B22O����e���4=CCޏ���??П/������.p*(	���>���D�>����$}N�K B4��������p"Aw?����?������)�s&�=�������������ߚ��ۃ����1��o��r���&� �B���@Pk��g}>�1U\>Ϳ��E@N1��oi�A<Ipz�����W�.����jxtJ� &׷lR�{�����_�����1�|�k��8�_����q��g��. Ed(�r���Ԉ��Eu"+�(DMJ��DWP �aEs #�]@��DWR����
.�u+�@]@��PP����.�Eu+�]@��TWP ���(��Eu(+�Q]B��R�A^k��Ϭ���|�t�o�ϣlct��{��������|lC	�!Bz�u]5��m��:ye�ٟ-��w��z0t�q=$��}G��K�:{}�l����v�v#6д>:f��k+K3U�T�;��x�Q�u�55Ś4n��=������xw/��h�~��w�c+�77[ѓU�ܖ�)�1nC=�j͚�]�F��.��*�ˢ\���g,ԦcQZ�3L���J5�b��0��a�b,h3��o�j�:����2,cO��;��w��H�]�	e ��q�^%�:S�<�z���Ԛ��98�W�}r�6��w���'�%�K�N�
u�e�1יK8�:Y]��N���˭燘G�Qa�A��찙B�u���J��U��x�Jt	J�M|,O$�|�2���J�C7��UhL^�0R�<�[�B��BG� �h0@f��u���ay����s�U`�I
�d2.��`ne���F�68E�F�6	V�5� ���c�2�S��I��ZJ�-�ugZ��:��G&��EɶcZ�צgJj���Ti�ƫ5q����&nq��X�k:��6�����j$��G�1)��}�߇�x�����|�\�! ��#3�|B"�I�G�YyTJ���}��Y�������1i�0�	����o��6x��Yw^a"��x=��{�^|D�of`�
�-:�h����mS�d]e��᳼����vGI*5Qj2��#*w�7�)fY�YZ:v�qޛ�c&��/�M��ݛ�*�q.���<��4����X$�eq��l�.�FQ��k���>_{�w��y�Wi�k�LO�ݺ��ݦ�'m�'nDo^�>7�$ ����k�C�ucp���x�ߴ�MI�9�i[{���Խ]��d#�����f�C@�������`�2�.�a�����3�,��-�����%"b@(J��J(J��(J,SF�7��R��g���/xi��A��ivMz��߭�;���o9�nU���4����S&��!��S55riU�d��ȸ�T�$�����N���Wi��cg@�v��h�̐��ٖd�Y��S)�{���,�y�f�����I,2�M5��wm݆��ь����2�FVK<���Z�]�f�L�."���QD��DItk�F�P�֊Ƭ:Ō��"��X��c)(J\F#!38�Fv2�'��+.���c�T�:pe<[nQ���[�8�/qL�-ȦVS�֌��V����5j\]o�/T♣*-�^4dլ�S�͊\`JL&K�FɘJ��6iU�Mbk#Ú�j�b��<k�Wo֥�O{�9Qj-�e#�ńŲ�gb:]� ?n �J\��fnr��̆c*�e�h҅=_$$ٽ��Ӡt=O%���8)�1&�t������(J��)��&��:�#,33���q�oq���eE��Gv���Jצ�K�<������)�zQ��Y�Y��M	�_,�K���rQ���N��w@�{�=z�zh@�!��%���^8
\XR��ǹ�;�qN��}�|�ű��Ř���b�G��1�1e���e��KK��k+Z��5���V�=e�W��[Y�nlN������O	N�a�}��%	BP�%;��uls�M�5[U�-�K�f4ڶj�X��[�n$�P�Ğ�ݻ��H��K�-S+��^��&VV.�=�gZ�k+3�y^o��K=�qMY2��e���j��X�,-F�L��樖�)��c�K�g�ws#J��^\,deMwZ�ɶLԲ���ܖ�&��5�!7���_:j5Z��d�\7Χ*-E��c�����˴���c	1b]�rrm�Y+=�.�'f�}��7��Y[�Y�;c�/;��۫9��1AI��Ѕ�6�h��h��ﯯ�8�.��bY�&7Be݈�6��Ф�5G��e��Δs�+;����V��s;�2¦2�����f���U`�ƥkKc%]b�/z�q嵇*eR�d��R�E&�4%	���g�>����^㧄��a)ż�*�06l!�;nq�ã"�vhX�7�_m�`�Y�c�0�QN���Mh��I1s&���UT��>J�BBS��N���N-�M���HؤG���ŋ�/��B���ugj�WǞ68R=C��h��)��7�ܳ�6.�[>�'X�HՋ�խr�j����/C<�U�N�B4,��f!a�u��w*ۼ��hX�w@��Ӕ�y�o3[�h�^n̛��5�߅�u�����Θ޼�����eUYy���u,̛K�Ī��7f���˘�."����o������rL��g�:���u��П���t4����C��88l ���6Fεku�P�Jq	��2f���l�2F7����3	JP��ѭ���XA�m^��a0r N��|���\�9ն2̬Ҙ�̧�qj�Պ�7T���B`�C$u�ׁE�8|E*�`5*^k��]��ǜc��=� �Ҟr���,b�icq�Vr�g� B"��!�a^����@��ݕ���{�1��෤uC ,')��X<|iP!+
�a{B���y���',���s����v3��Utݙz�{�d�5�e�z8�1�;ė��<���Y�B�-�{m�r8���O��s����v��*j�tj��ꗙ��4�WE���+A{N��j�{+�#�v�q��Li�r���.��9��m�f�*E��(Q��&w��Ƹ��8޴mq��
ȷ��;ɾ�Y.�n�$�{:���a���g3�wc��{�����.�6b��0=��=��x�V.�+�Mx_;g�@>ǝ��<�Ew��z�רXWӼ��%��,�<Y��M`�hM�_O��~y�O&�%�]���� �Áuk��vkG�ŷ}˻讎�X ������]>����'�A%cH\�7�]���#3�z���wk{��3��:c�Lj�ׇb3s���wc$�<��gl��tOW3y�.!gom����>I<-�7��up��Ƕ[ԕ�����g�RM��e�T 6FpgB|�|��P��q��J��Pxk��h]!��T-_��֭�T�l��)�"-g �y�V@ �Y&:�y@��!d���Vz���ɥ 	�_�p��{K����7�Ǯ��E.1����uml��2`��
��_*�Ʀ�$:���[f8�<�NfL^�j[��M��֛U�d��GU����j���e*����{�8s35Ӓ�]Y3n�#K���Λ��ڋQ�g��4���-�%/UK�1 |װ,��|ݯI����R^7���{ٞ/�;�c�e�L�u��-���k���7�˂�4.���E$��H/8����v�s���0[n�m�燴��胶m>���U���e��{�����?������ ?��/����dz:=�{�4{=�w���������=�������l�=��Ɵ��'�,��o������ 8����(���� �[A� ���@
P`8 p )�w�    Y@    ְ   �� ��(     ���G 0` b R��s��-YL� ���\-���6�UT�T�Y�V���mS�:9�X-��˗��=����T��-Gn��V����<�IE �i�8�����m&K�M�M.�h��T��V��ںwW $���  ���@H�@ -�) p���kh  �mk  l�  m�o ��m�^ r�  ���  �a���m���Z�Zlj�9�[u���J�^H� �tz7[V�m�mk� i͐�l �,׶��U�������a�nUU���� 2K)��H�.�m�W�k�\$�2��Vꚫir�-J�=R��yl�U��d	'�P U��gb�{�z2-��W\��%�������l� m�:��]m��Hd�ͨ펢_�g��mk��W�<��)@������dز6	�����"�6Ͷ�E��5v�u�;!�[F�sJ�@�����2��M������wG]l���l�n�`6�7kk�nq]����(w-g��d��@ �PRʰ��s@F�:m��)-UPpm��  d��$    �          j5��d���h�                                 p     ��   � 6�6�h �<  -�   �I�   h     m��&޵�            �� -[[ �        knE[@    @�x     �`     �^�7(ꪕ��uGhv�{u.��cӧ3ו�\�vv�-�8�]΅��r�olWR� �)�5�mN��IZ�S,�t�ܼ��J�7j�tΜͷ�~�ٱ��J�BٻH���j�J��S�L:G\��d��т�fŻG�m���㞣2����i\�m���P:+.�(��v����줡H�j��A �]�Uv㋇]"]��K^�%�fWd8�`y�tp��fM�=--B�U���m����m l �ە2 l��J�f�F�VqͶU�i.d	�Nz���j��/f��ô�um�86͔�B�)&���]���i�V���._���;vn^�x���P:�ڀ�mUs�( v6 �9k-��T��l�;��)<����]8���N&��F�H-�K5�F��a�W*�
�`�VڪWH�W��.�W0�J�6W�(��� �[uԚ�>VO�.� ]�Ѳ��YW�)X�Q�{f]��n���u������j��B�ay�i�
U���t�[mJ�tM%j���\YA!�uv{@:�`v<�F����4l�f]���$��V3��9V�)-��k�ҥ��.+��U��j`�ck�Lt�m��Z7I��RəV�ۭ�;80�:K���R�R��t푰�V(U�-�j8Z ګ��)wg�q@m�5�*���5Mي���k����h���V,�K���,p+,8Z�^:��病��-l�Ң�&��=c�V����lɭ��i��$�;rNj�J%J	N��2��[�v N�as��#�m���) mm��[t9B|� �@V�A��������u�*��A��j�6�M#m����苲�m��$[� 6�ʥ���dWAv����7hr��
pdӶ�;qu~�Wx@o���{嗫�eYV�j�j�C���f<�y��mًav��X�,��@�k��:�r�٫��e�%�Zl�UVں͌����歧���U.�n^`��v�z��6��t�nۥ��ȋ�f�U�P���Y�]���U���kn
�=P�da��.S��H[5�
N�Y@&�b#n�j�]�)���r֭�l�V�V���z����U��pq7Rg�̋�2�6MtٞwV��&��d$�F�5IwZY-U�4���jZ[��2���T�Q�v�Ymhf�;�v6�dj�umn"L�Ku(�具�T�����R�HL���Kv����k��ld.Ug�Z���	l�tV��k脝$�]j����6�m+�W��[��O.\���� t�7$�]Tn�u�Y�2�	XX˱�����^�Xwf� �l�D�;3�v��`j����W`蘠�.�mJ6�l�X!� v�KKY��Ϯ`�v��g�-�n	C�]�6t� .i�<vf8ݚճp:앳1��;a���
��vU�ʪV�xN�`�U��T�Y��^��N��s�`%gn^�Z�@f����m�sm�Cj��%�3��O]�f� u�s�E7E�)��6�s�5�'Pe����6ݞd<�4�l$�� �l�p � �`8(�T^�Z�h�mm4�Hi2��T��]J��u\JN!��mpm&�]sm� ���t��m�����ɼ�{M 6�`	.��[�uP^[G$��J�޺A�&�ۭ���β���jG�O8���\VԤ�ivkv�,`
U�4���ss�V��f�u\JՎ�5J���UV*I��i����A������"y*ڃŵ3��Ď���j2-+�6 J��.�ڪڶڍ
�u�J�ܬqN��s]��@h���[J<�i��� ���me��ZL^� 8�%���,v�j�U�J�@X���GP��A��UmQ<��m�`<7�x��{	 鰶ͤ�m��ڽY�zJ�v ��	�Ѫj�W`�U�|N�˃nAC;Wkn������c�P�8�٠5X�f�l-�l�@��������Mp�yN�"�[<!�9������ݎ���������:���_O�~Y�@Q �w����s��@}�������������A�v���P_����|�g���~���9p
Q>؅L��#D��$>�����!���Q��>��G�Gn��ܑ;�T"P�È��&	�H�Hy$6�xO!PM��VT4�H`�ʎ��,0R)ҥ�8����)ʈL!$C�!�y v�!PN�Hz%��C�Qw�D�C�i�&��4qdTV:�� y$ܜK[�M���*�ё:�m	"k��&��bE��dIa^��e���,�l�$!�6�9 S�]J�Јn��=Im
Z�*GRHz���'R5"c�������&	�<���'�$`���Q\�{)H<�Ob,�zH��Ae&5' ��Y4.�&b@���BBFA����(��$Cݟ��������D�J��=�|}bO�bJZ*Ã��)$�ĥ�A�q��	BR-BeFY��n-,��Z	BP�4	BP�%��Д$BP���
2�$��	�8��Rbq���`��JG�(�,JŇC�)K�����(JV�1�Á�\T`bB�)JH�(J����h)(*`b a���(J�@�>���3����h}@���w�M��l0�6� ){m�m���`q��Y��Z��Hsms�K�jM��l�s�@��U�U!J�q�� ���n�f݄�#����iԆh7OK���ûQ�SE�0�N�cV���k�(�v�.�f�㪃>,؋PS���n��	]6�� ��ѫeZ  &�&�      �	�[p�m	 $�� m�[�& m�9��������.q�`��҈��'V��e�3Cӹ���g\��okhn��Һ��4åJ��7��çmΉ;k�{&�d��ҡ�ΫJ��h�5Ѕ��ǵ)�rX��AL�y��{en3�3Ő��3b�cYnf�,���1=&m[��;�80@p�,Z[�����tF���1��r�n}`�D�pA���k�L���;s
tf�U���b������Y6������0p�!��x�v�r�0s���+���iqʱ��$)NM��F��u��Ͱ�͘1��4��Bi����J���,��m��N@�T e]�ɖ�U[^Q�S��\��3�ч��
b:ʳD0� Cf�]Y��6�`�9�J:� �T�4�jAq]gu��I���\��֮�q	v�n������w��������rH�=Hy>�`Ď�>�9C�@�t�ȟ�t��6�ɝ`���F��EC��]U���e�K�l�pH��_UUV(=K m�{;�hmЁ�Ql=�cg�T�Ǭg��wd���w;�8c�m�ͯI���>SV�J���wOV���iKu��i+�����̓�N��!ٔ�e��M�=�E��q��v��6�V-"q7��i��mӟ�T�Cy�Q�F�U�9�6Fw���!��Oܳ�Rf՛�＂=�A�^��zI�BiW��8zi{���?{��ȻMY/�]���{ګär�.���"�V��n�`�.��3�p���m��N�d٬��g:���8|G��8.��h�q�8��u�4��Ȅtj����`�i}��V�!m5^�����yV{ʹ���ػlM`��K�U��
�d��
:ѻ-f�EYު�ߚz>���}�zd��KH�tv'ے6�:�yen �X�Y �#y]��wu��K�A����i6�M*���He���yS���Yi�v^n�<q����+�u�^��.��1ì0ɳY� 3�@{ڇ�k�w�oȢ»�Ｋ��p�ֿ!�a>)++E�mzt�%Ōq��5�ez��[pجf�	�\���枏g}~����Y����v�6���ƺ��=�^�P�:
=hݖ��Y�*�� �$�0��,ζRһ�슻����(T�!�=��d&�o��My�V{ʳk����wds,,sє�F.5n��pn%ˣ�5�����N��ݞ�('b��si�%�f�b��U{�C��f�#~EJ��*�5�yW��Э�B�ht�|�N��yV{ʳ{�;b�m[���3�����*�<����3v�v�ͨ��q-%N|	)s�W���\����說ٷ:t(!�2������=�[��s����X���2�؊T�.1�c�Z�x��q�v��Q�.ur��#]���-�������k`Kfa����;�Ӥ�<��s.כ�YJ���[c�#H5�#s}y��.r�Y�(�5;gz�܈p���Y�[)h��Ｋ��8|i���G<&���m�KJ��=5'g�����Wb�4n����\�G=�^�a<��i�l�5��]�U{<�a�m�M��j[�c-�t3�YL����hz��	��^++��]�C�� I�^�4+l����|u�,�9Hj��-1Ria��9�M�H7�[e�~2�:��.�ռ>5��z���=��شF�B�<�Ov�dC4V�u��v����sP��^�f�Y�HYV��8�8S\ٮ\�T pܞ�%�V��Wp����<=����O=u��u�"�4n������CǞ��yD��s���V'�����d�!���>5��w�oȢ謭�*�j|k���GB��;M��<��^�{�T��}��} ��)�v똕w; �ƥ�/7V�Z���]��wO�w�CǞ�U@9��:�@�M�&��:���3����Rwj��{|���g�{�?{��Sh�SBP� ��9��T(Р 3�W���l��ѻw���;�<y�g�c�|�&���-��&��n����N%N��������n��C=`{0��%h�+��*�j����GAM�,;M��<�v�����<�{�^݂�j�6 7z�r*��Bs��-�6����g��X �=���,�X�%0�ہ�\v뗆*����v�6���j�f�u.! 8��2e�ݻ'=n�(x�K��{%��\��Um�ܠ�==��vnض������g:6��==�M�;��_����̵{Xf�`bc����ާwn��<�m��t�s@����7c��Ѱ-P��Z�ʛ6�_;��*�j,{�?z�e�Sh���s���`I�S�T��]��v]�ﮇ;�^�{<���~�;3wR�'�ouTȆKن�ߑE�Y^�*��X�w�{ݺT��X٩]"��Yx����8�L�Z��a,n]'�_P��{� �v*�l�]��j���WTWW{<���=��شDޚ��s���@g����l��H�W�ʻ��z�������6�mSU�ysP�U�yW$���~�j�[j6닜�lܝs$�F�p�f����w���*�yS9f��vf�{Uw�U����'8n���QtVT�U�ղ�O�;q�N�;�q<"es�[!����1Ic"�QE>q��c6�`
-�|��6�`Š���ż9����\c^ƺ�28�6Ȼiˮѫw��O;����a�%8��$��LSQ<QAC9�&x!�$wD�ùBQCB����R����̴ ��T܃��N3�pd���B�RF,�\�R��%�bΤ�:[e)V�C�����Xo��v7kI! ��)�}�+���j����t�Z�e�M��6\X���4D�K:r������1'�4��*%�s}뫯GŜ���vxH��
v��
��p�(t	�k�`�d|�'bx����I$��f�)�q�̧]�ʔ�w�9@җ]��Xֈ��gZ��P%|w�ԥ)�92�#I�|du)@4�N�T	��l�]�i�x�+��Ts�L�JR�s�@җ|w�)@�END)��MP�
�vBCRd&բ�[�e�]�����;p�Q�f�S�G[l[�ɬ�M��)<󼎥)K�9Δ�(|�̧�E��;�R��ɕ)JO\z�3޵gV���ü)z��t'�����r:��8�&T�)<�|��:$1)���k�A��8;�N��8$��_���\I��u)@�s�t�)IǞuѓ,��6�6��@���=y�(Ҕ���GR���gJP��>�@��dQ8 �@�ALM%UP� !	H� �����	P�%4IAAESIACP,��%���JR�s�c�u�F�ce)JO^���R����� z笂��9U��(��p`������!m���<�Z��Ki;9�Β_4+Op���.��:R���2:��7�9T�P&��B���'t]ݶ�i��B����#�w 1)�s�i�$��P&�ȘA��͞�+�V6ֶ��)Ju�r�)I�<du)J[��t�!E{���)���;cF2k5���i;﬎�iK~9Δ�({߼��(;$9�r�)I���֬�X����}�JR�z{�Ҕ�>g �F$��du)@��=y�<���s;b��xw�n�+���oGW\9��L>�㳣g���l�KUPF���r���r[�X�13���1�E�y��6X�1�7�k��vҤ�2�q=�����{9����ӹ⼑�Y4������m��[�F���\]�k,cwߒt���|'�Uh��i�+�x&2�t��jJb���s�?��t�GZ)��v�Uj�"�{�u)J\s��JRw댫�J߾Ӫ�hM��b�ü�HWP&�zd��B�@4� Je):﬎�)K�^��)[���E��bJ[�c�u�F�`�JR��;��R����J�BH��>q�WR��>dʔ�'��X�|3�i���)@t�)���:R���򺔥8�&T�i<󌎥)K��wm�-�meP&�*v!L�h���	�R����r:��-�~�t��Jwz
[?��lcJ��6Nz��5۪�9v�A��ܣ@o9|V��ƅt�ET��)I�;�u)J[��t�N�Yf]JP���GR����]�ɬ�M��)=z�#��x�d+�i)Ju��w�)JP��9JR�y�*{������ˣ�z՜��,l;�R�~�gJR�<��GP��	�O]dʔ�4>��������h��!�XO�h@ #��L�"���$ׁ&���&I��z.�L;��\$�D��
���=<�I=��2I��ɒO��A�]�O�z9��{CkU�����g;��3 ��)����}��g���������~߸:N��T��ʦد9ɚ����,�3�i��z�^��H�( M%)J�$�c��T^�ɚ��k��2�BP�J$�)b3~�7v�"ݴ�O��d��A��+����Q)�I���K�d�!���VMB5mk�8w��fP�덵��|�:�ۯ:�Y��gFq���w�C�$�`�d����'�$���2`�D �W�&I���b�h0�_���$�6��d����=�g����4�kX]B�X��-ے6�FI�%�ak��߫|�z��)�]�������~���餐�'$����n�n�L���WB��PD���d��|��P��v}�P�0��p���"Ow����
�y��d��ڐ^���8F6��I>�:u���z��:���3����>K+#���:şFs�6wޫ�^����IH����y�f~��@=��7��\gG;mveIl�]c�@tc�p��:Y`Y,�K|�5�7�ky�o\�y�Y�W<��^y���$�!�ګ�|�$���a�a^f5�O��4E
q]uƵU��gU^y�uہU�
&�U�}�e�h4
I��6I9���@�4�@�&o=u�U뼙�o.\�Sbѻ�	�
�ThPK���'�ɒ~�>�(���>l�7G�춛v�w�^y�uW���\��^o�U��gUny���i���;S-ve�5�H��LpZ �ڶ�\>�ۓ�zk�A��'1�ٹ1�+A��ڠ�jzu�c�c2Ɯ���]��=[��C�%�m��hSZ�,t��=[5��Y�]Y�x���m�Ѡ�Oku�]
������|����n92���u��gd�m���xP4EP|�p�v
a��x�I��'���^���y��1+����������Tcm����'w�I;����R�<�:��2g��dH�T�y��qg�9Ɯ�}��y�U��t]���Hwt��}�4�~��@?~��jU��u�m]B2�ʖ1��Uu�L�y�͒h
�@���ɒOg���0�k;�u�L���o�v���3��?|���mw�F�e��A�P��R��As[K�˪��߉:q0s�Š�(a'�ߛ$�n�I?}��$� �/Ǣke6-]��	'dL�
��	'|�$���26@�L�h�I�m�$�<�'�� 3#d��$�Ox�v
l���&����$�5�I䉒&�I<�7�l�,3v0�;$����d�&�I�A����?]�
�n�`R�57a�\[��.,��ҋEv�hx����%laip�.|�d����=�����6I}�|�L�w��߾O��@��__�aN6I�}�l
��B��ߌ��F�f.}�3E��W�(ЈdP1y�|ƪ�禍f��LZ�,a"���>�l�=�&I<�&I P��I�z>�e&m�����3��#�D�	
�s�ޏ� �?���O����]夭0Y�M�H͖Ș�1�3pw\��/� (�
 
 �:y}h�I�-�����d���;�d�}��=����1�w̽gz��&} 2)�R �5�]�Uz�>�Uo��u
�����>�ZɣV0mW���=���lB�~�2Ob����V�_8I�@|@G�d��D�<�I�(ȍ�SEP4�J,0��B����Uo�wf0�	���I�d�9�"L�l�:������m'�h���ƶ��l���¬Eٰ�}��-�:�¼�����"N�[$�(]P$�H�'�u��I�X�L�l(�uid��$� �_���N�]�8Iءd�y�L{D���'��3�i;n��@�{"d���&�M�P�,���6.��ݞcK����'�� ="�'/��m��uW�c�uϳî+ٶ2m������w�%�*�2�)��%MSI2AQ3-,�]��_��N�cz2M'V�ld�d*���L�C�%%����$�����q���K��&� d�����,��8voC�Qɠ�[:�YI���"+�y6&�e����*c�\�<�:�H��9�t��D�L�0,�8:�9�c's�`��f�B��1<��ք�f!a��	�b@��:�[a��A�]�4�Z�-%����֥I�QWg°n�u<���]��d��ٌb���9s�J�i��QaU��t�%�]5���x�eL��3i�*�`R���`��m�M�vPa���m�p6��$p�e�2��]\U�E���q��3���G��+�td�j�)L�-C���k�r�s�
�X���I�zbkS�@��^K���,��mt(���+4�ݵ��Y�RD�صʛ���Oj�cm�f	)cR<����^����I��  ��      �F���v� �� ��t` t��p � �l��u�}�I��X�<5۔�l:���g���qxC���:�Љ� ��^C8��e#'*�Q�i�l�v�flsҎ^ϖ�6��k��s`��p��f4:ч�M��"FWm-v��Ў#h��e0jw<�9��r��3���]���a6����l쨥�p��[��R��Ԏ���e�j`S�9��n�\�wU;X4��nZ��l&�1�Au�%.rJ�s���Yuۛ��ȭ��>�\���`�j�vzCѠ��y�Ol�It��ى��AҌ!0Eɲ333�㇭������i�77�~g��|�[�<���c�'�
�ZlCUR�uS�QT�KKoW 5�Ș�*�;K�۶� 9 ��eꉣ�����M�v܅-�ظ��U;82��ڭ��٦�Q�=��c�&�;=mZb�33�O���:N����GuS�N�w2(H^��}' ���
�T"�����Gٗf�J��̱�0��a�K�d���巜�vn����͋h�д��ib�öG@j���I�7;{ �[[\�gny�hL;���Zb́�[������]�6���l-�����Tm�[.^�nu=X2���6��9�������,u�x�;j��:KYwn�l펉#+$�F	��L��-�I���'�ZY$��4�	�~��$���~����\�'}gկj��0�����ꮽd�^�s�Uy든�,XL��O$L��A@�gcd�E$��}�ôѼ��p��DѢ�ߚ3W\��U����Ґ�*�1߾L�������%�$��$��P�(�:�ګ�<Ϊ�̙�������X�p=Y�X��v�KG`5�]
��t����	:vOS�Jlۮ�:I����'���=�I���}Ιx�V���$�ȟ�6�&�GH��+�Ier6�R��n�ˍ���iS	:0�I��fHGp��{'�
���3W�:֪߼�i^�b���뻰7vy�.g�"Ow[�R}'B����߲����QэZC	�� \���;�ŒN}�d�BQ��"O��ol��V�p���ŒNo�$� �2kd��}ᖅ��,�D�d3��N;ym�v�oJ/��x~ |�l�a2�8I;��d�j���ۯ��2��WŒO{>2�;M��p��2g��(P��]kUy�|�U��&I�wI�Ťӳc	2F�9޽8x
!H��
UD�*L
�H�B�bϞgUo�Lծ��9֬��qg}�Чj�dY_^m��W��y�O� P��3�~����;gj�<�j��
C��5W�z֪��}H���	�h��7M[\۩�nl.�3X��h��Uv�#B
ݞcK���"Ow[$Ψ~�d�}�`>��Q�Il�߿����{���$��$�� P�?oE��Z	:K�$|�,�s|��UUw��D���d�>Ӡ�,XM�g	@�}�d���&�L���G����aZ��V��G��M���'�I����UI	>~���߲<�P�M�͒e\��P��7�k3ۄ�H�L����vla&H�'�ZY$�L�؂$�	���i�v(X�	*�|��؂$ɭ�@9�/-�i;n�8I<�0I2kd�E$�J�A���$�A"��A{��'�B����2O:JE��d]�$�F�4(~�$���d���$�9@f����N�n\�Xv3�޲�Z����a+�x�ٰq-��檪�7<!~�*W���ɮ��6sև�U/ը.uՁ�àZ��-�;�(8Y�����b�	��1��Rٴ�en�jg,�1N4Se��S��5�;���vք��]�ݒ�d��eݢ�\ZT���d��\:l��}���d����=����~ߛ$����Te�nI��߲N��$�C�S|�$��6I����'��붓Ebx�M�y3W<s�^�Q���,�n}gժ�}zΪ��<��ь�Y�,P��B�H��#�]�֪��j�<Ϋl�� �@�	ϛ�~�O;֬�՜��G~_I<�&I�Agcd�=�&�mX�Y��1��S�n�OAg6��V-k:��V���m��Ǫ�v9< ���@��L������T���4j�:#��/5j�l�;�י2��Pt+�ï$�P�	<�L�
"�{������d]�$�>l�έ,���Ug�|�'~A��z����t�8oC��z��Ww�UǙ3HzPǮ}kT��O���2ܞ {��!�t���_�~��=�߄^���|?i�[Ҭ]��ͻYCW���3��g�m&��y��L�����<�B��t�{�� ~����G4��?}��Ԓu�O��=~��?~�O��~���6��z��vj����	K��C�X�x(eY �35�O��/*�-Z8H�{"d��&v6I�
$΃��d�<ė	2 �?���~��$����N�/��C�6ﷵ��.e�7��a�Lh�pnNU/��|��|�tR[<�����0����X� �3z>��-�����O��B�$��d�D�5��
UVL�}vm�,&m$���d��'ﵲL�Q$��#n�M���Wt �I��d�.� ����]P�M��&s��b�;60�$r�Y;~(�s"d�D��V��-F�l���Ԅՠ&ι�V�&���T)��1��ey�L�Wn�ũ�dA
���
O�y�L���;*�:��_�\�]�t���L����񞀕_@ȥ�^�.��E�V���s�ߐD��l���I.D�<��4Yh7��(#w�z�\c�5[w�u^�B�}��7��W�ZI���$�I��:���f���Z�p<膂��pɂ�B��H�2���o�;�3��s�y�ő=<Yn�)�m��h�3�Jb�)� �ch�-��f��x���v��	̽�{DN�r)q��3l�ǃ~����~c�5�lr'D@��@,���s�.`������y�Pmp9�p�0kW]�{=�ٮF\�n�����gH1�kI9�)[�8�O
�ri�X����$�3��FXL�8I;�$?s��,�p�O��P�]��)�b\$Ȃ� �@dﵲ����?g�wIgu���+K0���l��҉����2H�A\=[(&PW�@�D����>�"hQ���}މ�ݴ�j��I���{�"L�l��?�_���_��lrep�t��N�G`F>��|�?,�%�H�I��d�p�S'�n@��?}���,��/v���q��V6D�p6C��W{��U�( &s�Z�E���|�&\(�{�L�$�~���� �~��ң,�q�w��2OuI�$˅O2A�m&�y�	2 �$�L�.I2jdpZ���e������2�h��>|��U�SC�\-�d�b{�͒{zQ$���d�d�I�z&�PL�W8I�
�I��d�%�K��O��0�h�h�$�$��wB�W=F�(�{1:���a|htK�Yd�jw�9;ݱW�2]u�����Rޑ⃩����a�t2��4�VಣuQ�0EF�� Ȟf'>:��tV���z���#tZ�S.E�F��թ6V-�鑪��kvZ�i䧰�[���LR�T������:�I�lsgMS1KAD�l��������Q�z���=��@�W#��+�>'
�x��!;����D��D����S����G/�f�ٲd>���P�>�I�y�O��D��ڙ$��؛d�e�n�	<��OoJ$�52I��'���c�:C�.�əi�P�R礯k6��[GBN��O�	2�(�wu2I���vN}�d��޿�vņ�$����Ov�윑�L�I<�ݴ�M��\$�-_u�L�Q$ɩ�d�/X���e^$l��҉7}�S�I ` ���Q��\��4�,Em�3�&s�v6�`�e� �]��D�����PL�W8I��(�w��$�t�9#d���u l�J7k��И����T$+ffL�8uǀϿ̀{�Q'${�L�Q&p� �!��.L��9��&\(�d��<�(Mm�ɻ�$�F�'��	�S$�%�O��Z�E���|�&\(�wu2I��%��'nO_�ݻb�v�	'�&I,H�7x��V�E�����LA�7χ�5hD�h���2��7.ٵ4����XK��)�a.�|�wEUV�Yt(R��
�K;[��0�uA��+E�c��W8�`�5Gc��,�F��%'��T�0��Ǩ�q�7���˾+����*�mh����nn� Km���l���4V=an�X�P���:�E��j�����˼I��^5�O� �/�˲e�P�����r���Y��m<���p{�I2jd�TI�=[(&Q+�$˅N�P��I�$��3
a��V��Ed��{�"Hr:�~'��d�yw���AI��<9�Hƙ'�e4$��Λ�����Ք�iZ`��bͲٳx9"�檓UP��{:%��m�Żʝ�ʠ$PCqXɕ0�LRA2��iCCx$��Psʩ�m����$U��ES"9�6�ci7��}UB꾖3|���W�j�}��:�I�e`䊾�y��yW�{����|R�k�Y�\��/i���ih�`{��dJʝ��uT�Aȫ��S4Z��$U����D��E݃/�<�n�uJ���T�*�'�h�l�E��*�j�؅�:���Z�F�L[��ث{���"�M�z��W�$삮�(�֎;s�D��n7k�e�M	����'�w�d��D8s�m�Xշ��T�^<�*��؀���a[v�X;"�檝�����ke"Z���b��}Ut����r�t���v�j�W��V�P�dA�p�����v�7��[$�k��b�zk
�YMvd7�ҩ<�n��N�\��Mm�Ȼ��w5'b�:��4ZZ���5�;nj�:�ȕ>I�����ݬ��^����U�|�<�v�5m�U'��5TȪr*�x�:i;�Y6�*.����	�P�k3��ס�-ۻ^ $Ύ)e�gn#��{{\���>�m:-����J2���gYCB&�s,��*	�ZѴ4S�E��V텖�[3J�H�X��pk��\N�W�����Ro��g�:t�%����R+tnv���aИ5Y�n-ME�h��O�n���_s��C��Ml�]�VT�U��Y%�9{�3U��լ�ȫw�N�S"ǽ]�1%Ry�S"�P�<��]��~�6ˢ�}�w5VH�N��Zl�h��7d��:���CꍝWb�f�&S6��F�L5yS�Vn���b\T�!���ņ�evEڨ	��1
�%!J&��%Q�D@Dm����C��S<�U�Ͼ�K��,U��W{�z�P~�ʹ�ʦ|;gXI2�{�]�U�*��d<[)3h]�N�Y��N�;����������at�[
2�8w*�;z����4:��+Y]�V�P���D�zػ���iT�C{��EY"�9ڗf�t^	諹��ܪ�
� b�U'�z%��ZI��*v*��Ru	ة�CgAi���슷z��U2!�����D�l0Y6�l��٢����.����	�fv�ZO�O���d���vΰ�e�X'�DM�w"�:�x�Ml�͡w�;f�:��U���)��-Z���{ڄ�����
 P�ȸ�C�v.��9��I�/{��"��VxB{wi�}d	Պ9�t�hXv��͖�Hݶ��&
�+��}�n�j��T�C��6���L%yS�}T( 缫���Ͼ�F�	�n�WdU��9"�'"��x��yj�Z�RywUL��"�,�!$�7kȀ����w�}�r{6#�y6;Y�����
f2�b2(B�I��	�aa�e	��e�%BR�hhHB�[��K���:�!keH�\�+:ӗf#(�HyWVh�@sߗO�0��A��-�n�M6�[P@	 � �����l���C	�D�e�;��mm%pCXжv�l�fh�˳�kk�Wm#�h*z�R�9�W@e��v'ɰ�'���Ԝ��f۝��v�{.3�6�W0���֞\Ś��4�/kuum
!��Mlh2Ai��� t��(      � 8[@H$۶ ���  �q��	 	 e�n���׮�It�L@�"�6&�q����.���;�ٹ:9�z��x��]�vT���6ֶ^$���g�#h���')�ZbA�2��arVhk*)���<�#���*�a�T]8�lp����p�����oT�a���8�uH�AK�.9'��۞�´��j{ar,��@1�a\��U�b�Q 9���-9��9A6��Yֶ�d��q� ���$��!��kÀ���pj,q�;&L�k#��ZP����V��Յ*2]h��H���v�02�Z�s����q�;��N�P��st��,�k��]�3��A��t`U�up�]��4t1��H����2���[�-����������j��sj��S-���Upݨ{R9�kR*�N�2T��,i&�a�Jvp��Ƭ��ƶWįt��N�]�M$�z4���dd<���HG�<�z��d�������6��Ö��v��>kvNùцf+��n�v �A�j��p�P8�d��	���9Z�-lW���·��;s����u�ڶ��/�n�g��.'�z5]f��Fݫ��,����T���m)6�6����wt�R��,ew0�R���j�A�,Η55i�d��e �#r��U��^��9"�w�iL4�j�Vȫw�rES"� pN軱w�(�ZU��n�4�ϕw"�A��
&�vm�����[�*��*���	�E���yS�W7UI�9"����v���̔��͌�ڬ��$�$�I�m�6XL[v��E[�C�*��\�f��YO-b�<�]����p�&%21�S���;s�����j�,�!$˲�l�����*��d<[-�U�ʝ����N��{����i�լ��V�P䊦D3�Bnʱ��Ѷ�[��aa���-��i@�i�@�v.ز��Ry��dU;rv�(�eٷ��/�P�=ث�qW�u#�w�j-$ūʛsuUP� D*��`�]w��Ｚߞ��M�ݬU
#�|���9�ʾϐ�\��ye<KI�9�U2*䊾�>i6�����Me,P��l�a|�
M��M�aYl��.�蟿*�j�~��$�Y��lf�b����3�g������0�E�X��[�_�G��*��!0r�,������W�y�U2!�2����;w`��V�.ͼ�WsUN�Ru���{%Y_Y$���hދ��:��
��N�Zm��-�E���|��P�꯾�"����a0�k*z*��"��eɠ�w�S�X�O!��S"�H���3HI��"���3'P�=͖�*��N�\�U'P䊺�u�IDVSv�R�-Tj�7n��i���㶭�����i��T��]�]�i�ɧcr�N�;@m[]���ۂ�����I�����iy1�-c��sn)��k�N(�
��b�vƒ������ɼ\ˑ5���7Ktt���N��tb(|��nB�����k�����X,6�����l��i-����� &D=���"�S���$y��r*䊟</��˳oȫ���KwRu��IZ�@ݺ���wb�:�~��w반a���|�7P䊧b�:mիak�%���I���J�b�QI�i�����x�*�s��v*䊦\���a�x6E�LUP�4�ުr*��x"�m�U�ʞ����"�W���Za4��*��9"�؇��M�X�MWdC����\��}�'O���[�_֦h�����a���&�pe봤��i2�������UϾ]#�k����6�b��I��Dw�UϾC�|���}v��&v�EOuJ��Z����@��uΰ(� (WO"�N!̿{A�^�%���;���\�W 噤$�i^�U���"�"��-�n�mݰӴ�Gl\���ͻ3h�e����*��"�n�r|(U;�ʧ;���a5k+~�S�C�*�P�v�������s��MU�d龈QI�n��WwUrD���]�9;.�����++ވ| �G��\��9�ʳ�U��J��!�B4�>{Y�.w0,4l��a�wiݢão+dU��rE� ���;۟x]����߾C���b'� 9l�!$�J�l����$@d�g�Z�J7yS��P""��K�L4�wkȀ�����߾U�|�C��S��H!)�r��lf�� �L���ኑ
;gA�n����c�	3��W+["�����`3�¦i�R��͔�i���kV���W����!]4�v��,j�D{�v5ٍ�iCk����{<GR�.��
�����d;�I��Iy𑸞BMtյͺ�6I�-&N�"���pfʬݻvK�rD9�U;rD'�B�L�v�l����;"&��;gZi�&��@d�rE\硲��6�l��C�*��s�&��sN��;"�U;���;�d�w���m�դ�;p�=mge����璌����)��e�|�*��w�H���%��%yS�: ��
� Ufߐu�U8&�h�k�@su�W$A�΂n�(�E`"���!;8o�Re۵�� 9���@rD;�C�Wb�^����0k�K�;��:��i��V��M#m2W+�P��G$C�*�&�kU��o�@su�W$C��4]���K ���9(_�0Ѡk�	��2x��-МD9���´�\Rg*Y�I��1*�f�q�7��fXʜcSZM���Ɔ�3'HtI:�/B6IH�e��@��ܡ� �$EƱ��97�&�b""�ťMk4�&���*��d�ij^��{1��CBx8A;^�t*/ +Р#A�E7@����.�������4��-+��su	؀�?���an�D;�@rD2E\�ӲR��un��KB�6�f\��\�0�Qnd�t�,��=�C$U��9�&�2�ݼd_@�*��!�ډ���ZЊ)6]��z*��j� ��:�H�L�����$BPC ����ЋZ��x$�n��U��>=F�V���[4�l�lY��5�Ι�mS7����ݬdA�UrD���;fi	&]�x9"�n�y܈d=-����h��9"ES�n�a��6�I�@9rD2v��[*�5�s�y<���g���ǜ�1£,wIА�~?}�
��K��f���b0�Q�(c9Mq��6[u�fj���`���\���.�eP0ִus�� ��ee4;<k�;g�O.�pk�����!��!��.��׋S����q�q0;aS���n�M�@q����bt��N�t�'�a�'��X��Bu�aڈ����vRmV�e�.֎MU��j@�}��>v�6�%e}���H��{����6�	"�����b��_��`�%7k �=�S�	5 ����	&ZW��*]�'"g��o�'���c=A�O�%Ʋ�] ���;mۻ4��@�ʞ�wu� �U�	�e��-Z�$C��!b��L	;��]���8�q�=d�����f�ڼ� �UN�$����"�M�k$U��j$A��k����W���2EO�W0�z�х�lڶ�% ���q��;NEnB�v��e;��b�x$���_ k�������ӵ�w�9�*�~C� F|;_�$�j�~�W{�� �P /�h"8&������wP"E^���Xj�j�	"y�9NE������bY�ѕ*i��j�[��]���eY�iK&͈>�Ȅ��rm���d���E]�&�'"��i#m2VT؆�'"EY�![v�o����Oc����i��vL��Zwz���/h��`b��r!&�2	d�m�7~�.@�� �<&�~��|^��7e�t�۱v-����*�5��D�C�:ذ�7�6!���AȽ@�ú���Ds�� ��*������+eZ����9���b��s���D+l��rE]�&�'"��`�� �Q���),hȅ�~=����[�&4�l4���B9�5;F��1�t�@�f�h�+1�V����GP��kvy��9w=�à�T�.V���&�<;��jOZƭ5�dt��B�u[*���DQBλf��#�����
�ɧh%��2�u�m�Á[y��S�t�h�pjo(a��C-���T�[uD'U=���q,����[��r!'g$:]6�ʓUnjqT�_ *�צ}�m&-�6����!��S�U8G,�!$W����:�j}���8$G[�x>?}�y���~��w���@/����֠XK�ݫ�J5�ж,%,�ae��K�@njuT�A��v"Vʲ�;�����*���*s�vq�UɿZ��B��k�yWw�}��'"�:5�H�L+��O ��	���\����찞	5P��$�:���;��|���^�id7>U���L�h�6�-�31��m'e�Y^3R�U'P��	�9ޔ�M^	5|�j}���� �t}�>lXB��G�ު2���7F��ʪ�ϗ�����U��K��75	8�N�;ޫ��U�x�C��Ru	8���"��Yd�$ވ�Q�G��*����-&��LYE[d��MU��q2 �zv�6�
�������u�>C︫9��K�ٻa<jsV�:�Ρ���H�ݬv!��RuP��X�Ro �9�w�6�J�zj��
� ����� >��������i�)3��nٍ�P�%���K����z�t%�o ��n�2!'{�n��ݰ�X$��'I�'{�v"Vʳo ��wx�N�';-�Ӳ�	5Ww�I�Xg"��i#m0�*O!��Ȅ�Uq+�.��IM7N�m�9,9q��������-6
Z����D1�1�Qj5�(B�(lR���"��&Q5�PD�-,�g;��Ƀ�b���k4\�/NZ�8�].iqW5��7�LY��S��/3H���/~v�l��q���j-��]�0e�uxyb�r���\m[c�'A���l�p� ��A#��8��U!��N냎��Rڪ�BJX�0���*�dj���5*��,qT���	<rj-2��8�tݰ���8_n�L���1�ƒµCUT3�g�Iu������՛�-�Y�$؝�\��K�H-66� zt��     � ��`$m�p�� �� [�  �ěZ�u��c��mR9SX�a+Xk+��1K%Ҁyvn��в���2�<���$$�b�[Vl�M/b9�&�@��-�UY�R7d�m�#[��	��JŖ�T�r�E�՞ϘKmd(蜷k7<���l���3�OD������î��u���9�y�qd����j�l���$C��<�om��k���D�4�v�z^̻gg�Qg���T�!��F2�F���V��ձd0Q�{V��7e3���V&(V���t���(��SJ�u`��[m��κX��"�=8�;�5L�-s,`Z��X4�s�Pg	�W��E�ogL��Zuj���'�`��ͩ=�����G�k����$�z9��Bb�R���%�l@�cK$tǲf�C
s�S֎4�����'ޓ�:H�O��5�t�>	�wI:w�;�t���s*�HF��w��*T�F��;	G`��� ]K�r����1��R��
ݶu;{jK���v۬�D�P<���$&�df�4c�eYL�D�[n�7^#Y��s��<'E�K�ɫ^b��8���Kk��N�|%��m��4��!�2��ܙ���0�M7ve�M�m����}�=�Z�5A���N�v�H��I�I�AȮ���v�����I���"Du,Y��"�@9���8&�*ݰ�j�'I��UWG�@�D|V��:I�\;��F�M�R�-+�ҶU�|�|�w��ߪ�}�P�~��!ӷk�jt)� :� 1�HI�����M"�b�*H��C�����:U(�6�x$��'�P＇L�z����k ��!��Rjq ��عq�m�ͶJ�Z�פ�z/-���Ӂ�;Y��i�j��BN �g	#�b��E[�@9���\t[vö�I�������}��?����䭕f�T�{��o�����9!Gim�k$U��$��	+�h�n�d�-0��hh}��7	�/�WE3m����+*H���"�d*�d]��	"
F{�g�*��C���ڴ�n��}�> ��}�|9�:[l6���߾u�y��(`����
���o��:�	��" =�03��n}C�?M��\�KH68;!9Ƹ�&��+u��5��m`� �ERj9�v%�f���9"��缫＇�j9��B(�Mk$U��$���g$�F�e^�T�����|���t�Q�m��#�Pr*�P�����M���d�L^96zwes�%k�Rn�M�<��[��ܛUUV���)K0m ��&�nx��Tut�A{f�'79�Rۨl�Қk���001&L2�Ћ-�a�=l�#)e4���6����݌T�r� ����ϑ|������~j�㉱�9���/7m�%"��.ê��.�|���n�N}���}���1��@g~�>-�M`��*��jȾ��:,ϑh�W�|��� �U+�n�v�m�D�T�C� ����w|�õnɷ�s�{���'���.�n��ﬁ�X��Bu��=BZ<M�^�Ln��k$U��I�"$�4��ʼ{�gn��p�c	eFW}�1��7���E�S�Z���Y$Y:����2�${�w�'ɦ��_���4�_3wl��� �W��@��_}��m��&����!��^���P�'E�m��kdU��N�4�0r	�T��{���\�i���>�S�蘐xՒq�=��}=��ޚr!�*�	��]�[e`��i*�P���vVѶ�H�n�f��VT��)$h)��D��Pr$&DN��,�I��`��l����}ߐ��H-^�-�U�I��8�H��z�х��fմSV���.�:e3E�����:`�Ϛ�mۼ���d��(���0�����X~�w���l�{��ƹ>�6ݰ�w��E[��@��o�>�s���U�ly_}�u �C(
�B���ʚ;��L����w��T�C�d�/�0J��l��v�WA�*��PKV����w�?��C7UI�'b'b�n�I�v^ȫ��'b�'�zV�#m2�*MC���C$T�+��Fͱo�@n��T�A�;�bv���$�3��N!;p�ڪ ~��?�]�[hJ��1	�4w`b]x�P�\�^�3B�0�f�UT��X-�.]�I�eݲ�=UY���.��ڹ�4�ɠ[��A��sB��Īr�C�~9M��X�9Y����X�*�j7ZЎ0��(n:�2-ձK@e}��]p�2�\�ջ�����m�O|��|�����OE��a6^��ʷx����Rqs�Ϣ�vlyRj��N!�/�@��~�Yb�-��o�|k}�3�*��I���+h��k�P��Rq	؀�H�Z�Rh�x;"����jN!���Z$�a
m�n�O�h���VXQ՛#A�ai�yRj�$�"D>J��1����'<�H��0��ġ��Yir�JT��azu�i�����3��E,�f�&���Rq	؀�A�m�Se�슷x���Rqs�Ϣ�vlyRjU
��ﺆ}� (O���~}����,�Q�vqe���٘qJ�+-f�re���>Vkw�?�U'���vVѶ��ɨ=�Rq	؇ �w�&���~�W<�q��41"IHґwԛ���U�6ֲ�1�<���D:��[����N��t��%[�n#.��hZر�����܂����N(� �DU���wd�ֹ|�yֳƆ�:Hu�D��EH|I ���D�$,)� ���q����u������kB6�*�5W{���"��WU(�ݲ^T�U��$�8��,}�i���d��b�+}������M[�31�ݬ�yi��P��T�U2 �=���E6^	<���S"�8��{f5v�ڥxh&���Rq	:�v�,Ze5m�N�]�!'P��(�J �#��)`S$��۽�[Y�D�6�a�-���MCw��⩑|����4D����ml.Z��ܛ�d���57	�gb���V��?s�Ru�L��MʓW�U7�U9�}�Y���|�ݲ^T�U��$�:�MۻX���U��U��5S�T�Cm�v]��*��S�S�	g+ 4LS�U�$�a	V���d��T�*QI�d���Hl F)�lw�}���s�ݼ�NRQivU%�G0�rE�r�K@�pg^ټ�uo���A�G�vT8ۮ�<Or�'X��ە'\rhRٳ���x�l�i��l�Z��	��^����F��y.Lgi�Q�A��Xf��m�k��#�{��캋ot���y|ݴ�)3���ٙ���lt�V1�볝N�C&�ݻT���ک�}�K�Sݷf�)���"�w��2yWf��N�����mW$CwP��5S�W9�Z�Rh��In��2EY�rK(��Mʒ*}�S"j�!��a^���
�����|�3gq]�ug%>ZM�d�v u	:�
 >��}��{�cڱ�[c;e��3�:hS����Ѫ��T�_P�D}�C��	;/�E]�U�|�ȇ89g�]��+��@��W��O���,Ze2�T�T��I�R|�����ˉ��M[\���8+0��0�EvG-�J/5\�ު�~ Pu�>U�ϗ��@�e%�ＫwUL����Tgw�-Z�F�e]�}���u@P�U~�	:��+���wl���@���7�}�U}����v��l<���"ު��S"��7-!r�
۷ъ�Q�s��#{O����7h�vR&M�O*��S"�"��\�ST�*H��<�>����Ϗ���L��9SuVwP��&��ٶA�/4!��7z�MA�TEF���B�QW9�]�
vRX;"����z�︼/o�z����L]����:�;;�:���-�*H���ND2E\�]T�7v�yS�S $������m���W$C;���S�T�=@�����vE[���K
�s��Gl���MVW�D/v�ȇ$U�
�$����1����-kE�\M�i(�V&���ɍ�8�z�mӔL��4�u*m��n �����·n-�nб�&Q�<�1X�m���5&�;J[��bur���x�\[f7��:�N�8�' �'&�s�#�qa̯9��t�V��@�ZA���!m�N�l�8M�v����M;6�m�����O��>�iy��"�!o�䋾��U3P���=i����*��2]9�=.�Zi3w�$C��t�C�!����(�ݰ^2]>��*�P�0���X�n�;h�3�%Ÿ:	ƫsFy��v�;�Ǌ�`6üN�!��7�B�&:~���|�KB)��o�,��4*�b��\�A�ԃ2]=�g9g�]����";�>@�|�~�3㺘)��X4�����I�{�6�ݼn�$y��N!�%Ӕ'U�k]�شӴ���^��b��x�;Y�%oE;),"���8d��P��Ϭw��W�-&n���p�n��H��,��1���7}���= J�C
��Cdj�Q��	�jo�i����x�r�üYu�$y�T�C��jN�RЊh���W7P�k�!��A�4XI Š�m��-�K�i鴺W^�M�n�j�%el����S�z*�C�n��ۼ.�uH��!��j�iۼf�D9�C�*���!߯�Ns�v�N�K��wP�C��$ P7wt3��
�4�z�z�l���D7��Ԛ�$U��퐔L�6����n��ݺe2ū��dY��	�wm�����C�/�PDg�!�>�,��L;x�}�^=��d��zpޒ��m���*{�r\5&���2+��@���s��pȐ�w�M���v����9"�"�Z�G���z�(r���&4&I3=�D�Xյ��$�,Ǒ�����IP,�(dW��K�3�HdfF�r:�/e�Q���v�ɋ�"-י(��4nI����ؔ�k�quq]�K;ŬɑU3"�M]�O( {��tA������k�}�=�_/���kD6���m@8-��9�lKM��`M��M��`�<̹4�<��9K�5mUQ2���Px��씠�Y*����J�p�=�=���pL�핖�G�[;6��S砕�"��ce;m�K���t#��B�ݎ�=9�Ք���m�H�M�m� �ɤ`     @ �`$6�$��` ��[wm�  � �wJV��Z�kE��d�lٗ��Ƭ��]����d���� ��+��K;[����p%<�5����w9��??�k�>=\6�M�;Wb!v��Μi�ٻF���\�{OX�G%�Rv���Q�,�e:pkt.X#�U:�3/m�\�;p\'r2�sܷh�Y���X���1Q��
5s9E]��Ԍg�$v�.�Ȣ3�;	ڋ<�K�pm�����`�c��X��-�
�a�ǁ2݃Ms�$��k�ث&��r�Ԣ�.��Gk.��n'����,�Aƍ��|���֔���|13J@��&�٤�]hіa�r�Yr��@�������$\�SH�[sZ�Q�]j���h�JIa�,3���r�V����I�P�p�ʁ�,!�\CYv	g{*�89:㩎��I��<-�x�~&���P�Da�f��:��{!��!�&HH�;�Ͼ�|PWf�B�Y�cPl�r���GM�vݭ��ڕ9&�	28�kmoY0���#�*���	X�	u��IM;����I�lan���5\�$N���KX򕮋�ѕ�#�N�"���1Y�26�Lj]SV�t��t��,(�ip]s��
E9�xz��6��ݐ��m�V�n��f��wU?D9.y"ڻH�d��͑�o��5&���{E�J��soMI�rEY��ʰ�6[7�e�]�C�*r!�Ӻ��	0��5$C����r\5�����hYd乸�E9����o�_>�19�l��v�@�t�v�=�ʞ���5&��xL��a�rD� +�{zjN*�� Q~;�Ke��^W���n�D��9�0�V�N��#�R�����S��<C�/�g>�y�$�X7�>��I�O^Bz�\���e��5����r�EqZ�V#�=�ŶJ��soM5�H�3�YVF�f�l�k��N�NE����e��0�m���2s�9<#����R������`�vA���2m�;��7�-����EOu�I�>!&�A]�rD/;�	5	ث��tOt;�[V�607��t��uv�ໜ\�i�S,7j�vD�;�@���;�~�#j�Nݬ|b��
;�U�|�}���-E+	;&�	諹�`�#Ru��@��m��H���Ԛ�u�M�U@C#�0�bk ����xΝ��*�a�_�| ���ϻ���޿}���W�֤�Z����%*�]K2Tg����Sf.�����O�k�m􋵴�k�D�����Rj���I�F�b��:��U��&Xm+��/���U2!�t�V��o0�'�w5S�	/����������q�)�DpmH�+�ͱt�϶xܗj\�tUUn��@����g�kA{T�Z�#5��nWqv�7��h�f-����Fkg��k��,�+��l��^�)ac8<\�rm����cN}r6����ø�;�l�Z�4\v�N��Lt�p��l%a'd��;���$��>�P����>D�++�����ԝBdU��,�
"-��C=u��̸���7�R�-��;�"��ȇ�
��۩��/m0�5������Ԛ�N�- �m���]0�6*	ݎ�KѸz�'6͋WvY(0m��W$C�{u&�2*�D�Pl7n�C=r����yȩȃ�h�j�']I��P��>C��n�>�j"ͧf�}��ug.��3���:�vݛ��}B���ݺ��!��U��JOr��ݚC[5Q݁��n��3�;F����T�O���u��$�"�N�Kh��o��!��"���դZL+M`�ʞ�UUt ,)L�$,+	(�a6]��\�A��>aR��H�NmԚ�����uh(&[�x!���$�"'M}���v�y �z���0<tI1Wj�-�֝3�����D3uS��
c�]g>�y"ӳvV���B˩5S��V��n�"{�Rj"��	��b"�+�@}}u����U����=���w_}}�ND!�u�@��ؿ���a�b��c�m�Z�O��t
7h�a�ȶ�V����*{��?mԚ�a�>aVW$C�v�MAȫ��AA2ݻ��[��䎳"!�u4�qeԑ��Ȅ3n�H�"ӳvV��_nz���X|�ewe@�&�$���?M���i��%5�'C��ڻRt�X�l���a0���UUZ��=J�q ݧ�m�����z:g8��%.f�ʻ�V���Ya�t��=\V+(�]M�aLh��աtĸA
�Υ�0�ѝ�f.�p�����wI�t�Rx[����a��jzbt�v�n����㞶�[J�l�m���Pӻu;r*y7�D[eg2]n�5VH��^�l0�x���A�Ud�C6�=��-��x9"��B�S���}	6�����ݺ��9w��_��m�$�dh��ғ�d���ZNb�1�L;a$�A2ݻ���:��V{�d�U�i�d�˩�� �C-��Y"Ϳ�����6E�f�^�����n�b�Ԭd;l��vD4��N�&���Q�XM�,�|�>�V}����g<��'3�*�qnE�B��開��|��<�k�|�������$B�^�����j�H���B�S���BM��WdP���49{��M�\irt��L�Db(0Wy�Jt��Z,\�BPA&�����m�x��Td%p1��n�!���F���ơ�;��$i��Ұ̇Mn�"B�72��q�&C(`33�tso�N%�0��Qi�QcOY�g$g)�!��29�$�L��L��c#�@�x��A�f��8&a`��8�t=WM��a���wR�Y3W����n{��D���� ^�N��=��c�"l$�G����P���<��ٚ�H�E^g���Aȫ$A�iW��i��.����$B�{��w~0`��me��z�-��q�u'�ڑ��;K8�1���䊳��3o�#��}��`���o+�|��۩؃�S�	����+2]w���VH�ӻ��6���n��Ԍ�`Èp� `I�C�� J'w|t�s�p�n��6�V����Vn�;p��C�89��y��OB�p�Ӳv�����vf�\�!*�c���i﷦���d���D��E�*�O\5��"���m^�l��jz!���D'ny"Ј6�7n�vEY�Bv�5�Ԭ��w���ޚ�P� 94�M����)���a�6�5�4u��΃5Wm�v������R�EK� Pyçn)���T'U�g�����N6s�"�l{&�8]�h7E�CVx�q���g���r�Nx�kC��i�l>i:� G�v���w;�	�m�h�����n���)�9�^g������9h�	ۆ���H�����T���a��k���guS�	ۇ� ,l�K�6�V���ک��o�Rj�$�h��"��v!�*���N���ou�VH�=�V:U�Lm�`��\�<�
��v�;5YV��l��jz!���D'n�N�F�����vE�S��@�}�=8��b�D�vٻ��wuW�B����}�s�M��J�7�������ERst�a��-`DuS�	5�,Z��O�՗Z�b�m��-�?���_1�)r�j�s5]�{��s�柿jMC��&�@��������W=�3[);�M�� 7t+� n�<�S���Gn�-���zD�"��+�����A�ѱo>�S�BM@O���n��o�\~+�ػ4�I+�r��t�����+�z(���H�wP�"�s���1���D�Pr*�I�V�,6k RF3��ȇ��9'M�&��w�:�򩺫@�khd��#{��VW$CwPjE^�&]�;w���wib�s��,3�`[��d
˚&�I�Vo 7u"�"��ݦ[7o � �U9�PӣB �hط��*{����~C�����v�x<m��Cv�k����U�x}F�Jڻ�=p�/�u�"�� P���!m'vKۊö���YNLf6�զ8�u�7:���/$��nxV(lp�;&���'=` ��>��v�R��P���<tv��k�'O+�])�f�Ex�e���.�f�(�3�-]͍�Ћ������J��,̽$�7W&�[���d���֎E���!2�|y�
�ńy����U�!;p�$���i0����#;�M�jwP���F�D��Ȇ����C$U��3[)i���/�{|�}���3�j;v��v񚞈<�u�N�^�5|�7K�4m�����pX��CfR��B�ZW��������v*�P�a�J�v�y\�%�UUѕA�^U��C>�"9��Q��V��T�U��d����Ѫ�1a�������!���ʾ�ʹ'n��I�m<�W�+��_oʾ��?�C��i�5VTnك.̮84r^��m���cS�O��"���W',�l�ͫ7�OE��dU�+9�5�M�yx�OD3u	C����71Tȫ2j�h�j����EOuT�C�  ~��w���%z��A��}��UI�d��M}%^�I�]�	)�Y����dƭ�ӝ���ia+a]�OE]�C$T�U&���ņ^b�"��Ȫv/�;>ۿX���M�߾L��U�~U�9�a�F�
��H�{���;��]@���ʬY1���ZɆ �"�SK76���a8�+�sS��2���R�7�=wu�S�ᮛ
Y;y ��K:}��x蒡+m#l;m�զ�ǍT��r*���$W�MY/dT�UN�Rj�j&���ɼ�H����P䊽���p%l+�UTd�V��g�!�>�W�xhW�A�,U��| �[&W>�ϾU������ �S�GԔ�������?�`D�`�( 'g��`�����H]�I�\d����la���9�Y2]㋍��6���I!i(�Re�jI�"��IeH�p@�.'�%� fA�
- �$WЀ�AS��H��JTr@
b@iJS�@��B�� ��Ωv�@T|�S�#H�lIh����2n��-�	䪘�F�V�4��@�!@%+@<B��
Esu�I��$��$G) wb�����R !�]�FSiP-�*�:�`UiDB�����d��y����Qݎ����$�9��oG�~+�YKa�,�P�"P���!T�\��3�������:�����a�:�_�;���ƣ|��q����8�D� �d�OҘ�Γ�A��]��m��~E�n�է���O��i�i��~���c�?��z��=BC�'�0q�td��~c�_��g�E�]��c����o��O�M���u��|0~���ov|;�����|�?�y^��������<������������}ݒ	�-�'���}���?W�[��G�����ߡ��a���Ⱥ ������o�G���f;�z���OУ���$�A�������ӈ�������R�}�W�����qh:ӣ<���9�6:�a�&�o��c_���Lpc��Cw�_����4���D���n=������Q{�rDr���������}7ݞ/��\a�g޲?����@QW����}���p�UBTI�p �
H��*$���
@�
J#
$
� �*0
H
@ʉ�� ��)�K ��
J� � ʉ
�
HH)@))"&8QI�THH!	� !��BU��H $BVBX,,���"�R��BU!$A��E���,,IaD�PXTI,,AaI
�EQAQB��,-P�BY	X	I		BaHQdE�RQDT�a`J�$�Y$��	��$ I`!$XY,EXQa�!E�*B���QH,(�E�
��QAaAaRQQ`�aUJ$���!�%���QRY$Q`��P�QdK
E��XX,!�*
� @�HH� B$�B����,����I I!,�!(@2�!��*�Y	
B�@02�0��!,�$!! g�¨fQi@�B$"@�� I
(R�X�����,0 �J�I ),���
J�
D
$H)*���@�]����s�{,s$:�~��߼�A�xz�y��&q�����~���>)���.A���iɺ|~���}����0|N�r@`�>>�ݿ�׀����kO�����'��p�G����{���D�c���9������O���B��8d~o�ɴ��#�Ԙ���>��o䏍��~��o?n������؝j�lm��VJ�����ƻT�?W�������r��&�������c����|�����_m��~�����f����
v�d�A��槫-�a�Ϥ}?V?�k�~����?=�������l�`�}�?���c�mf�,};�@�S�	~�}�$��>��J��p}�r)���:�����m�Ly(|~:� �}pn�\lTL��N&}��~�ч.�l�A�?�Ҷ?:�%{�}��?O�$�C���90@xv&ìU%��+UK�b�#��7Bu'R��q5\��F��#]O�rO��s��9G�Y ��Bɦ�aO��:���������K��k���o�H$�~���?g�?����~���Ƿ��- ��>���_ۿ�����?q�?�s����O���A��_��f�_��_�3�>����?Ii��6XO���/�߶��������F��A ����z�E��y�'���ڡj����G��~[�aOd�@&�z�O�k'��{�^>���O_��=����-�t?�dq~π{����ϛ�:	!�'���1�~�w����1��޷
�.5����1��ˉ��'a'������t��1��t?��p5�>��xtr'���c'������P�9�X���{$XŊ�����y���N,`{:7��O���Շ�s�c��w�h�l����ì����>l����_��;hC�??�������#*����!���G�&�>��(}����;q���!�}�uT�/���g��n"nh��������x㻬/1��ݸ����'�}���?>����{(��I��z��G��]��BA�L