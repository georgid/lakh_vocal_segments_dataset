BZh91AY&SYÓS1e߀ryg����������`�  �
��   � �4 T �  � @��y�  ��!��!�	UH
�T�P )
�TT��   n
 �@�n�{:c-v����ˣ\Y���8%�g���@�N Hz�$:�C ��OA�(
p�R����{�>��G�GŐ`V@4}�}��/=L�Z�p lvç@Ǹ�xU�����]����0_oM��8�����  (� x{��ﳾܴ�n�����y��:m��{�_u�M�_ 6�ۯ^��`}/}�v���{�^�|�>����n���]׶�{�6�(�� ����|��Ե�#^����<ܜ��wMۇ���ݺ�w| 1݋mp^�i��)���)�i�i�r;���(( U �����3M�ní:|�G:lk�ϧv:�@	鮝t�	��=�Ϻ�ܾ����v�5���_x9i��ϓ^��+�              4�Di�J�FF	��0�&L 0  щ2���)	�2L	��4�A�z�TB�F#CM�LFA�FM Ob�P(J�        ?B���SP�44`�d`L�LF �"B�И!�z�4h �i�Hا�����|���>�Ϳ���M EP��XQ��ߥDT�����S�8*"��~����?�4*h�_����������o����n�o����|��������c��?���0��:�����f����߮|��BI >�*�⪊W2�S�#��Õ%T�v��ۥP��ȉ�y��x�h��>\��vWe+��݉�]��*�����T���N�G<����~~����~�N������u���u�	��&D2(	�@L�d  ��P" �� &E2(	�@L�dA$@ ��Ȁ&A2	� L�d@ ��Ƞ&A2	�@L�dC ��� &A2	� L�d@ �Pr	�@K�dP"��Ƞ&A2(	��"���&@A2 	��d@O� &����j��# ��s��*�d��q���o��I��&�½����QA�]JL�SL�J�5Q�e��ĸt�(=�T�:.&%M!Q����*BLB�h�WP�;���j�Rn��V��%����C�����рV����R�Q��
*� ����X�i�Koqv�B����!��SE�(�M��Pl*!U$!mV&�q�*�
�G�a��Tȅ
��G��a3Ԣd�2���jÖc�NA�-[F�.���#̱o*�����(�h�au*@�a�,C*�D�F�R�tY��x��f3Lc1�JƳI�����u�IH�F�e&�e�PjD*�XK�t��𰩆�V{���#�+�`|���76������PYq,�.	 �	"�	!�ԩW*�\���21.�)*�P$$c5T$�iP0{�A��F�Kq2UB7
��Wt����;2m
���$�H��A���@,�Zkf��ʣ���z�u�THG�I�wW	*���f�6ȕ�q����D:�2����g&�ү�E�Z%U!�
L��B�ǋR��.Qk��dJN��&�XYɰ%P�j�(��RM]����P*%A%Q��TA�����*-E��dJ�rT(d�P A�IPMU	"�4��d(p�a �	 RH n�IZ�R������5U\����V�B��*M7�a��iR��5 ��ʪ%�NK���+�+��7��%h-q���bB�ʡ#�) �) �w�|�ӓT�Qr!�@��$�H$�T��	 �	 �	"�	PMA7�$�U�y
nB\�$�U�BH$�L��	%,*TbT(e��F�B��Jm�27�5/,�s4.�h��N�K���J#�A�3�tg	K�_&���Bd*�2A&�XW&f�=��u�Y
���R%A$Kd�Q�Q)(���\��Q�5
l� Y.5�)P�O;(0	VJ�f��B�14�����U�haQ����BH�4oz�l52��@*�G!�2�E��*	!@TZj!TA$M�\�d!r�
$�R�k2f�����;eP��I$%Y�%@,��
��cpi�V��T��F -ĺh��uL/!��.ap�K��\l�$�TZ��*��r����n�fY�C!q�\*tMK˭+%fn^:u����D��d�B��I�CVԁw����&J���G*������e���neM!PI �Ph*-5���R埽�s��s����=�ߗ�뱼�$�URH�Z%A!�E���F\J��
���*5����,����r�F��	"P���)��S�(��Z")ªR�n�6�|L�xv̆��R�V�;r�'!tEUBD�7!U@e�
*��12�{um��5�h�)
�DA$(
�l��K�D*�B�\
e�#�,�a�NU%%A$*A�$�MA$:�$*6���˲L,ַU��¹f�����8jd*�l�ǨQ�z	��.��a�9�s�RS���*t��juR�o�f�'Fd6f� �{�O}g0��w�hݽ3�[�p�q�d�d���%E*'\:3��RL24�ơ�cpI
�e��u���tr�H_ye���^��$�H%TB�#�Ģ<�k�P�	���²��.8�M���d�I%WmH��yV�ܺ�jnJ"��ل+mˉ�v]\hmM*%R6�lTr=�����h�g.�az��l%���qe���1�sN�]TO����Q(l��w��I$����Ql*]^��9&���:�A5t�$�TZ*�
*��4\�\
�]�C���3��\������ĸ�N�C��m&J����l�\R�"bT�Z�u��jHd$�;�P.%`j:�v�\
�Q�(%��!�Sr�h�����KÐ���n)"��Ƈ.�M!Q�74�C�(jR��XXl��*���	�A*	 ���e%�G����T�ˮow�Yp�Z5��dh���f��5��4w�0�o�� VUɲ�btʹ�.��a%�.�$%q-*��d�I�K�T��	 �) sFC,��Bu�*Dk9��R�uK.�%H�����R����U3�WD/
2t�Hp{ܣヂ�Fo��Y��C��e膮��p�6��;ʃ���WaP�/�h�XK������P�
�Ŭ�|���Z�t�XM�$��H� F�
7Ui%��������B�������)�@���R�P�*	)
�m�F�.����s��ow3P�{ꛗF:�Ż�h�(
��F��]�g+.�����vK�o}k0�Z-�uE]G(�@$�U]����gE��;$���N�P(j	�ԉP08K��˅��CE��BG���
.��e޺aD��QVx����*N����<<�[�Rj�����72�z��59�	�Pp���(�B�T!U{VrpI�$�H��I�Z�of�5$���
���4�ˇM�ʒˎ��C�S���6B�E�K������IK�L�tH�K��w-�Md!J�}Bn�,bi�n	�Qn�bsmj%�T�9|�P�Xm�/���³�����Ұ�4j��	Pq�2�	Q)�p
��%K	.��"M�4�ȔcsF��p�e2�M^	�%�<������\��ʤ.	�:���B������w����E�9pI�7:r	 �	 ���z�S��Zj�K�UJ"I��km�-+���\�M1�%L$�VKu����Tn5Y��utj�@���p��:����U�԰��E�Q.	������A$�&���J�H��j	pK�\���J�T�Q���]n��um������SS#.3[�U�,�3D	�ڢ]݅l��Z%f�\���rH���a��-5(m��D�ԣ=��o�W%��]�QZ��d���ژ�J�q�U�bPԁGRt���Ǿ��V�F���Äe��d��w
�K�W��*	�S��'9]��|���B�XE���IP.%JB�� ���.I���R&�̼�����N�rY�t=���r��@,�IL�����@9`�d� U�?_[�n�����p��l?�w���������ݽ˟ݏG�Y�z���bW�z�9���e%�V�"�/�w3MgIVg�t�~vwŚ����+������?W�������a�ϙ��(3��oS�������OuW׸����}e�Q�3Fr���̺��ˡQk�Μ�;�6��(G��t��c��Ze�h����IH�Z �g�1��f���믰��j���e����1��!ڏk���F�J��R%�HR�4MW\��յ��d�dA���U�RZ*���*�[m  �[d  I�p     � ^�P	�� d   � J            �      ��@
P`8 p (0 8��  �J �`   3��    �`���\       ��           �$       ����    �            �           l  �{��5�ۖ�6�RI0u�!Ō���zڔ���î���Jʪ%7QU ��V��7�8��1YBB˸��;ajݬb���][F�pmJrm���� ))�n�ۉ��3�l�����I� [m���eUyW�%��Tթ
�`�`۶�f�[dm%m����a!ǆ� @R�ԫR�P!r�c5�X`  	�f��  j�a�H�B،��Zޅ������ �im�[�/J  [Vm�   � m�j����RZ���h���h��]n�˭a��   ����f�f2	6i�[z@m�V�8��.�u�o�[Ml�м���k�1m�� ��[VkvvK�C�|>��ߏ��  �g8Z(g���u�p�����K<���`�Ԧ2��ԧ�6�q��ہ̩*�+�G��ݵR�I�Ii6��E��&��v�m����@��/[���  [@[v�鴂�.��mm $A� ��m 8$����ݻ��̭R�J���PH8@� �7nbY@%��j]�e�����i�RԎWbZ�T  m��!��j���� k.]�_-t� ��HJ��U[*�s`-���J&����UV��K����Z��OcB[m�i��`Ӗ@Xf� 6�.����!�`��ZU���
��*���ҲDK�[V��m�{f�ʹ��݅�ܲ+c� �z�۶Ŵ�nB��Qm��F�u�=Np<[Aa��/Iv��@[S��ݪU�C�Y�UR��KU0u*�Ut8�j�%���T�6�,�k%��`	M�<��Ӯ*Ȱ�Mmmu^�2�c-l�/����U-e�1  6�i(�kQ؛��f��`��	6ݛ`�K�rC��P)��'{�#[�[dm�]��U���T9j�vn. Hm&��Xm"I  �6�	9'�� �6��6ͷ�r�K��UUR�r�[]m3k�5��Zci-��`-�x��� ��Cu�n��մ�t9���l��ְX^J�n���   E�K.W	ک���bK�N�V��Y[e�i�1�l��Zچ+���ȃm&$d-��CZ��U�V��V��@n�m�2I4�@-��Hm�]��e@X ���%u�T�-��z��ڶ ��`��5J�S���*�V�@�UPM�LsZ͗��/=6Hsm�7m�mW�	E  -��lM�	� V� j� nN�Gm� Z��˲K0p�` 2 f���Z6�z��hu�`	l )@6[��m��5� �	Х6�`��MT��J��U�*ʵUV�ݼ�@ekv�E�\�޵��­T���k��]��ļ��  m���-�u�WR��倪��U�vh :νe���$ۮ���[�&m� ���c�6��mZF�9m	8$�\   ݚm#i�M�6݀��86Ͱm�!T
�ڮ�	U��v�ـ�5�l6��h$8����5AKR��c"ˠ��hI$O#m����|��8�4&�fE���K�h��V�K�4���&vj��Pj�
�U.�s���  H/GH� �d�F���{��H�r�� � �  ��z��@ 6�ÀM�%@]��z����_��YI�m&Ͷ�m��@[@�m��m�   �` &�l��X h)@ m�m��l :    ��a�8m���ŵ�[��W�7m��ݝ� �`۶qm�-�[ >m�i�����-��� �� t� d�lC[�����mm��`m�L��hH	dP�kn
��B�U+���0�R��F�[\m�؁  k �t&�*yF �j�I�QΛ�Z�Wes�WRU�W
Z�ҭ��Ԫ�C�J���Y	�j��������ݑ@�RȂ����)�Wf�T��bFE��mf[q�������f&�Y٫�:kL���}g;v����ִ�HH����a�m��  � K-��kkj�e+6�h �Ԁi��   ��v�[�l�l\�V� [@[T���ʵS/F�J�:w
9�� Cm�mnZ��[��>}Y� �]���'T�ҝ��Y�]�3p5�n�6�e�ޝ�8�$�U�W+UWU[�   <-���  sm���6  6�/-�2mRm$���>f�.eX
y�IU�P�v$9�`9f�m��i7�QԫZE��M:�UYV�43j�]Rم� �Wh���l�K�X�K��$  ��  �ӤZ��  	��Y!���q���Q�Iհ�md�Ul�]0܌�ˑ!��C���3ј�G[)�uA�難�Yk���h[�S�~�8{R�*l�G_�ɒ��"���6�U~?�~V���9�'���;�u������g쿗�
�߻�=�_����ø~s�������t�?|AS�}~xC�|�߇�����_�}��S�q��� ��D�� ��Dƍ��� I�!�6���:5�^��
W��thw�a"@� �	�`BD$aD� @�	�UG�j�!�[R(�(.	 �@C���d:T5� b0Ua�: �RD
AP���(�$��H�t�G`*E 1TN�BX�,PCH�J\"ǈ�Q��$c$��b�H�`�*�J%�t�Q`��z�B�t�AC� ��W���D{T^���ؘ��P,^`�j'hȈ3�Ihpy�=�Tx�J"	 � ! 6��U��i�	B/� �1�:{T8��\K$E;Xi�@pT�b!i
Pt�F�pZ�`/5�
0�+�]*&��(�A�pK����,O����QE#$�a/����k��4��D�{D*��O�ʃ��
� 2H�,�#"H ȢH(�"2 H��*��H ��
�0��!"�HI! ) �2(�I#3��L��}a�K���.��c�Չ�v�-��sÕmE�vY:��9�GR�:P���`   p (0ll�@�� -�����    ��uҫv������f�g��<HR�`t�e�e�k>�v�b�YFyZ�(q�w� �M��W����Ai��[&`@ j�ː�8ba��ѱ[�M�K�w]t� �e������D�Wh��r�n� 'D�*�Z��t���h�@֦��W+��jD�U��Ƨ�h$�pcQ,p�vೃ�rSR8���I1����]���F��m�����d�)-��ۥv	��].��S�`wVYė��l@cz9l��Ō�qc�t%-f�m�f��`�Z�e�32�m5��*d�4�ZҖ@�ɚV���q�3*9ڥs��EN�A�57[]�YhMѧVX�w*����p�hx�C��,��+.���3U]/.�J�N�S)-+�`,�MV�Y{h6yv'��3�@9y#cʠ7u����v�B���c�j�୮Bv�����V�vg�������ey3�=���t��h��rVq�#����QWj�Znqs�Z6��#�MX����i���
����/ݶ��������9��G{�F���� ��@����{�	���ڠ�J��SH
��P��u��"�ڼa[m��m�s���kn$.�S����!fi9-�l�n�i��R�0�uX�͔�9�본�-����6vO=�>�a�l���-D�R�rs����1\vv�&�j A��8궈���p&��!��c_��{����¸���;���"�p;vl�Cb����³��sJ�?,]��y�r$�d����l��;�:�J�8ֻ"MD�&k�z��i�:c�ˮ�ȢD���{�Pَ�.�wk�t�R$�g:a�i�N�c���{��Q	
0mHӪ��&���g�/F��֗"C��h��;�:�J�\齩%F�R��;�RA;U����t��Y�^y�*�a6k�V���W��v+Er	��/k�]N����N�]Ѹ	6HƱ�����c���r�����B�����]���ɦ54�OhNF�cr4��BL�N�c|Ӫ�V;:�t��H�5;�<o+�uӺX�RL���W�k�Qb�����5����Cm��%�D�*��}���S!�^�m��e_�k�U}�� 3�����-�QXY�=,j��t��1mI���.0�l�ṣ߿�*�5��W���v|o��������^z��t����k�7&��;��ٽ*�V�*�4���l�Y.��=���_i��ʊ@�k������U�w/&\zs��]N����w��T��"q�ゞ^��eGE��X�T8�q$�g�Ʀ�N��]��tޛ����)"�u�ɵ��;�a�{���������c���v�]�]d���7����r��_?��ύ����K ��R���2u&��%P�ѵ��E����@A�rym! M���J���)�h�TC�O������63�.dv���j8�����6��.�m'Uay�q<�·�ʜnNg��;b��Ά�zo���gq@��QP˺�\�َw�Q*VdAM���s��}���&��0�`,q�����zjۥ�j��6��mZ5�=;u&��M.����(�v^ut�U�����r�/*�Ĥlp��{�鯟�?��z���)&IB�W���WLw�u�zn�F㤤��]J�َ�o��}�߿�� A��A�}=�Ǟ���4�is�{��WDM�ֺ�b�ͼwk�u��Cq128c��/`T
F%Y��KD0�����;��z�!�(��cSn�WLw�u+�7&��;���[1���X|��IjS5���U]�&/�-��VZFB�mEv�Ǟ�h���Z� Hp�
&������x�vu���`w����vJ������C!�Rj����@�ٯ��N��Ƈ�'�`�m���H~�e��-#�ߏ��U��;:��]⦙$*��<ok���;߿����|~�n�����K���݅�\6�.�<a�L�h��cSn�WLw�u��xs �d�k��M���v�ݮ�:ky��ALֺ�c���v��׎�ulJ(ӄf;�<ok�u�����U�C���6o���8�V56�ut�{��Wt���mJnbA�N$����,��z`���4�ZS@���� ����j�������e����� �|yT�Q��X�i2D��{Ǎ�c���W@�{���ʉHG��W!s�8e�j=��vJVڴ��u��َ�o��u�m�))��I���<���WM��{g\�vմ{T�Rwܻ?��;.��w�m��ڸ�ۉ��-��.Sv��^ѫ[�e+�mD;�L�h�1�u�=W"��VW-�ܐ�F�+rbm;��Gjs�%�潸�h.��׻����}�Zy�N�@�x9�X�Si�e�L��e��n�������SH?�}��K-����X�52 �_z���-�}�=R�C.����Cm��%�GU͈g��UM4�}㬶E�p{����[��	�	�.�q��i��p\hۛ�/*��]^8.��w[,r:������t���O���������-�Y_|r�xTURx��v�ut���R����$cX��ml�[x��뢌jS5����6�Wv��z7�eulJ(ӄf;�<ok�u:�c��#`��4�U$BqD��)eMY��u��:n;���G}��-���מ���{�}�!�ڐ�i4	m��� ����j���*�M<�a�Y���+��ȇ�A	�64�=1�=S�h!Im��(��JEE!B��J$��B E##�(�E�Q��l�vBlL�@�K���IH�T35�l4���ӗDB��o�7��XB!�b�(҄���qSe�u��0z��͛U�:�F9�j�����Ъ��@,�� �-�ECN�Ѿ�D�ք:�u�ʵ$RD���r"�����.�fdҒ# ���H�몵$D�^X�RE5��1I�|�y�Wuu����k,w�I�jH��ǚ��QIߗ��$RA�άr#"���*�o��MƬ����`䅞�`�q'��{ݷ��'���"�E7��1I�|�Odf��);�I�4o���\�ˬ�z�dS����$RAﾭr)"�ΪԑI�yc�=0j)�z�W��+.�&\ڒ) �ז9�E']U�"��z�Ȥ�k��b�) ��<�wWW�U�^�w��%y�Z�)"u��r)"���1I�C�>$h��^��ٮA�7c�I��]�2y�$RD�Z�R@"�]X/�u`�r�{ן�̘1Wc�P)���'W'Xf��"^7�(�������H�<�&)"�]�c�I����'���Ȥ�n�uR]�W32i�}z��!q
�u�ڒ) ��,r)"������n��d���3U���RE<���9��r)"�����H>yՎE$S^u+��YYXKҒ) ��,r :����H>yՎE$Sή��I$L�ߓ̻�ʬ�z�dS�_��II�;��R@}wv�H����"�#�Nw�n�ӷ�n?���Fk���U\�H��[p͗M�t���6�I�֑ڝ��p�q�x�q��%��n�e�Xv�Ckl&7v����-�8�]wn,앫��{n����'s��s� �]kv�%?����U��7��H�6B8��H�J�g:h��h�୔�����5�M3WS�9����6����o{�^wc�I�uV��H���@dS^_��I}�<�wWW�U�k,w�I�h{B��'\�� 2)�W�b�) ���ȧ��Uvu2�ɆfV��Iμ�Ȥ�k��b�) ��,r)"�ΪԑIG~r���3.���;�ȧ<�&)"�\��"�)<�I�<ߖ9�MW���]�W32iI�|��\�H�#]�V��H����"�)�W�b� ��E�RU��)u��e�]�4��td;]-�ہ��|�|?=����e'�U�"�7ՎE$S^_� �$�E$]z�Ȥ��EvV�++.UiI�=u��#=���%N��CQN�z����>���"�)=uV�ju(�L��sJT���G@& cL�A"�|��"�)=uV��Ȟo�\1@fվ	Ep���� ��ŕ��w{,裈ZYo@i��$6��p7��Q	
0.�7e�mŋ=`]S��ja(�B1Ĕ�d
�\�g���ݾwL���k[\$�Q5��vOURA�[��`{^��l�qSL� �[��t3N���g�n��@5o���|���ȉ/E�R^�`s}����Խ�8��]��#��<| ^��$_��-��ӊ��\��7&�4ڨ9_fˊ$H,������� ����2��r fվ$��8Fd�n s��z� ͻ ��:(�Bz3�.�z�fݐ�n�|�u�E$Y�r�>�n�nCb���D���5T))�S�{��B�c����܀;�C,�D8����\]s9y�I
�F*C�	bdT�$�@.�� s��y� ͻ Qu�|���i�օ�ΒN�W� @d�=TI�L�$���D ��z�k-GbY���x�C��\ �Sd׏FډTրߟ�����a�c^׳ 5��Ԕq����� 9���܀fݐ	�Z�j�S���
����[�W*U\�۫�њM�x�G��)��-3��zM6�:tmc��5�k���!�8���n��� v���?\��c���n.�(�;����;[.�M���HH;QqE��:��e��O���00��秺{륒X�Ɗn��Y�v�#�m�p�a�q��N�G��q07�H|�@ݸPj�8�B2I@�\��� .��_Wok���j&��7n�����V=���� ^ǎ&���$2�y� ��r�v@.��u�m9��3@i���@3n�{� �Q���VͰ7XmPI�r���C�J0	
B����qF%�/� �� /v��03�Wj4�J�A9��2�v�OI% ��3����ʈZe5� 3�o�(�N����&{�G�� ן��`p�d��Te#֘\�۲��n��7P��RE�/� ��
�n _��U���J&�IԠT��Q�|��k����s��0�r�b�$�ڙq��?����TA�z@4�^+����I�{�s�H;���� ��"E�߹Y�әʏ@���y!�UV�u��v����F��Y���k ww Nq@�8|Ld5e�ډRZ�Wj�U+���c�Lg��5�$�FS�HD^&9ݗ��Ǯy��f܁D�B�1Ț��\$��y� ʻP���q�N��^�.�y�e]�w� վq��d"�,�{� �� ��������䨚��h�� ;�8|L3U��T�X+B����j�u54�"��]@3�Ġ����w��b�(�6�����dJn����エF�C�i�&cNg*= ]������ .��݂�e��CY�r��(w����&����F�-h�� ;�8|L���Wȅ$c�5����&��V���0���2���$��Ips�d�Ku�I��W�O�˴I����q�E�2��C�Si��Κ<z)Pi����P �E��*@�d� k{,�R���R5� �F$�dy}�-�l:�U�nBF�l�H�d
��Ѫ5�� � �'#�SH������*P��
w �CG#ě�L֊�	``2�YDJB9hA$���6Ul���MK��D��tdA�0#�cg2�_��z��Q�RQ�Q�W\�n��r���#d��&J���̐n�l%M�    � �p �mp[B�)�   -��ll  �  �gE�O'j�8k�:����g��KS�=9��e6d�p���c���@vq7km�k$��mڒ���{mj7C���mNR�0m���/�u��L��n���zv�#��𝸴���ͤ��G6��ܙ�kP��]�*K]	�WN�qp�lZ���X.ya۰4��T��]
.�a����A<m����;q�)��%,]���ٯ'�scd<�H��˶�<��8ⶴ�R���F��Y�s�Nh-r���>%��7�VG{slt9��ÇvsqH��J�
c��*ʻDF`[:�^`[x�۵�˫�8Nf(�*4��&�������̮.�J��-Y�WM@���VF�g��W\�]�C��n�I8-��Zꪇ:[!��3L�z���!�p6؎']+��l�V��W���km`]���#δ�i����/j%|r0�+nU�q�}�w}������,�9�H�p�S`���J���*��X8��N\�m��I*��m��c�$��=��U�Y��h
�P�F���n�)���R�Th�"����p!� 8zE!I��DGC`��
����좭��X��m����@�u`uk%�s�9;0k$�I�l�u�B	�M��x�z_Z������ �S5�nϨ�î۷eni�&��C�#dۭ��s˷9��8�	�� ۮy7�݌�}:��k
ocF��\.;qS8���{޽ރ~ �
JV�6+�4b�*��[��ڤ�'���:�d"�,��_���'���y/m03W�NJ���ր����A�� /��y� .�j����c�d� s��Qy� ʻP�6�rf4�q���v��$*�@�]��3�̃QȆ������ .���05��X
B:r�= =e���yu��R%��v�(��M�5Ig@m]�����`^nB�ͫ�B�1Ț��\�*�cq@�Q)��ާ9'�W$�7�$�y�g�����+��PN��^�+�L��^�|p-���#!�d(�܀es� ]��(�&��%D�Mk@m]����P��y� 4t���YnF��[no<4���muq�]i||�}��#�揶������&�窫Td/y@/|��^LƜ�Tz ���� ʻP���.d�D5�/w \↩�1����)�z�i������{L(�h����_'��ݸ�&��6�|�RF9]��``���r,�� ������4�R9Pt㔜���u�f�s2�T�խ���'Zk/@ič�HUڔw� ���B2I@�܅W8��%|N��v��9*2(��6�j w�����I~�I|uD��*jBH*��| @�ת�'ޔIvꉱ@1L�� �r� �s.Esݥ�훤�ɘ�v�o<p�� .���~nv�͊ɑ+1��L�ks\q708�ɱ[$҂����q@�6T�V�:���(�%��v�;� /��y��-i+�B�28�@.��8���W W� ��Epv��/A�c
����d+�P0�K{�u�E$Y�r ��Tjw� {� ��UU�1���-Z��H�c�Ɠ�I�Gն�Xl��D�ݍ�R]ˇ6w;�;vN|AW=�[u�.eN�Ā!���||~�f���a��9�����cX�cZ;>��5xۉ��қA�[.�kIՆ#\�F2B=���0�Ld�ncYl�^vk��Ϥ�d���hn.y����"rTMD��W�� �ՌW�UY�Ծ����l�MEM�r,�}�\=�P��Lk���(���Grf4�LǠ���y!�1S�V$��� >���A�|���d*�X��iw� {�p.��K�L���6(�%�[^�� �$�^n@;����5U	�WR�&��uv�^�bIQ�*���4a�%�D)#%8ր=�p�L��}+�2����Q]��u���ֱ֝�g��rrv@2�j _x��X�1�U6qw�S�FB)"�w� ��ʼV1N���p֘��|NJ���ր��� �x��0��^פK����Tۧ"��� ��_*(wi������Psk�ρ6ӈ�	�*ٌ���f!l-�
�Kr�i�3�1�2f= ]��� �+���B��u�5��A��CY���UWՇ�i�}�\ ��������c�RZ��`��9Z�1U*�`k7 �\�B�14�UUEL���u0=�H��%~L���A:����&�U�k� �`�� ϶�*!,Y���F�9���n��pN�b(�S�h1���S�FB)"�� � ����t�پ'%F�mk@i��V*������Ɂ�~����L�����nE�(��8�&D�Hv��Gts&cNd�zab�L�Ns�D�ܢ~�� BDA$�H	`��"�����^I:�$��%��JP�ߤ � �ۀZ��{��[�.�z�Z�C���Lt܈��$p�x�gI�8�%��{ɀo�p/�rh5|HRF&�@.�������\�i� wZ��;j	և��-X��y!�1I�`�J�z�A��r
�ߤ � �ۀUU��f���MDִv���(V0/7 J�UF0cT�1  `�P4$$�B��Q �^�46��q�m��m�y#����I�e�u�b��3*'sq�M��ԧm�����]���yH=�7[����[m����'d]�ӫV������ I,tJq�gN��l;vծKI�c;�Jt%��T��
v�N�\���*۰m�d�Tt62Ýk�.��Q���R�~�T�q�I����Y�mp`{?Hv��Gts&cNd�z��� ��@\����$����Oon^v�BQ�|u��F���z@q: ����`L�{�j�փ�UV+cO� ���>_/�c�}銪�>��w����M,�}�\k��r ]�u��(@!��Q�H�(���[g����X�~?�v�{���=5�#���� � ��D��k�.�A��r]�7[�Ҫ�
QBEJI�:H+U�d�P��.倩� ��=0A�9����\���1U�k�<o��D�G� ]��q��UURV�03�H�\=I�̫�u�Z�E=�*�������]ސ>K���~��3s&r�$�^��"�{ @D"A�}ޤd�� �����,,���@�TF�S��\���:#n'v�q�����4�� 9��=�:�c�DA �,��I���*���8Of[�� �@���:ڢO'�i��K�׸���M,�]ۀmpbH�UZ�R��BD  H��6'W��(T�Ui&���� @�Fuc�QA"�ȪB*$�� F �222Cd�A!*PF�B��e8�b��$b) �
 �Q�-qL�b��y�WFS�eFo�T� �޵��M+�#���0���!M�ð�I
�tu��E�����2���kLkD����tu�N���k���=��K�c�p��-B%��PCJ�`���E�*z� Q�)��   ŻTI:�~�A+�4S�/A�ت_��a�w� {Ʌb���V)}� ھ�Pn(��B�{� s��]��-X���#i+M�N�)>՞F[\<�l��j �9T.@b��&��R�R�+�$�(�o�r����*�W�+��� �����R,�}������<V0�q�s&[Ref=j��$ �L�z�q��F�P�V]��&I<��;R)�u�����K�g	�qF�Ik@i�V+|�Z��.��V1Z�^�He9Q��BJ�D�[�٤Vȵ�c�n7�����YҤ�lM,�}�����>�@�����mA:����P���0�8�v]:�qD�2F�� �>��=����x�p��Q�@�`�ՌkJv�V���	�@.��6����0)xH
�	@���AX�I�I����B$"1q�`s�+euew�a2�*NN�m�����'FӖ�仐��mάݔݻ�R<j��SZݮX����-RT�mۯh�i٦��e�A��ݻ���m�pn7'g[*�r:�s]ձ��������g[Z��v���3��������w��r����N���Z�M�s�Cٶ����T	J�n���̷��L��ɘ��]�d ݭ�E�\��q��F�P����`q0�8��U���uG�z48��`�L|�yx`N܀j��ۍ��VLD~KmQ''�E7QM���ҵMBʵ�@ �y�mF�Q��w�����Tf��P	���9�iN+t��=e�k����Q���  <ho>��S(�������W�*�	!$��B@	"B(ĄH2! ��X����Q<��e��ݙ�����R�;��{I<����^�ookyέ�� ]��G[C���dڴ�U����춂�
�����s���on������H�%U5c��>�b|��Q�ڣ���+U�0>!�n2u$�A��Ǟc\�\n.ũ3!���Ww*�
 "�����I�e�"������E@U	����ջ(b8�}{ʇ
��Tܝj�j���p �*��Ub �mG������2R�d"Kʓ�B�wr�<��T�K�l��{�.����[����T�k�H��� �A9&qwo�I����}���x���aj���<�w !�D�'�y���X�j38��Q[���wҒ�I�����   ������^�ep2MR��-��o4�d�IREq�� p �	 g��y��ӫ���BE�Sq5I8�s��m9ؽ�T�O3���s%Y��[�Y���<݈��`
 ���p���jR�mFgn��/�� � `@ >���F�)����������z���$�F�T�Uq@0"j3�B�Q����v��V����@n� 0`�!%�oL ߻���MR��H���8��j݅WO9E}sX���En�y��W]�w,�赜txɩ��b��V�x�v�Vn��ռ�2#���>�3]��WoZ��\�x%Քs{q�HDG"-nɂ�������7�f�KA���s;o�+&��$+6�K[%��tl��8�m/�%���������@�����^JJ�2f��I��w�V� 0@�=~�)*H�W�ΡZ�m��zv��(Z�C���}�C��_�h�  ~��/���(�SR�\q�A 3�Pߔ7�7�'(T��Ok������;�9�u��& ҷF�۶�N����]ܫw�1���jrH�5"�J���pDLA!�Ey}(��o.�y��m�,��Қ��J=�B��}~ ��~Q�ڣ��'�b3IR�c�|���7q���͸Ѵ�6r��]ܪMAȪ{�w~�6���J����Q�hjy^,9��˾���˸~�"��AȀ���ۍ[��#���U��dU'*y6�A�L�S��nr�TbM4
�J�pؽmO<կy	�����%�����}��2r��a�+e�H'������D3'���U�j0��6c&�홈[p�N�E���o����xn�
�(���~Q���^Fi*T�q�H���Q��""���RU)�7��P�P����ɢ����c� @{����wf{{YDڢD�3۞�y����2�J��h<�=��o�1���W��ֽ�����*JJTR'R��7::��qn��g�3{l���e��H��!' $�>˗�Rv�)�5q��" � �{�@7�)�o�H�jEJJ�{u@��  1�m�����&U�*�+��D?|м�m � A＀޹8���J�)���| �g�7�:�?��t � =���
)�e�Ȣ)u�t���D�\�wfE�o���Ks��ѣ�gC5�z���d���d��\�Z7�Oݙ���a�E벋 �%��^T�� Y�p\�Y69�fH6�`�u��`   � 2 R� 'B� 6� ٵ�l     �6in��\�@qr�튌�H2�m:Bѱ �G���*�)��Y@j��a|�(=��uP:8��ܾj��"3��V��۪ �d��t6L�)yW-Ǒ֬��κ��*����BQ��!˽�	�l0)ҁ#ٱӒ��LMǶnM�C���zv;\��ڸ�U1cţOKe�8�&�&x9;d�����M&��ce�iMB����G�dN�:9���.v�=�5Ӣ�S��2J�n�糼��sx���$�-�n
Ӹ�ۅT�s֕j��+Ғfj��v�P\��KZ�=����nx�B[��X���j��[ ���/���%��l���� �ӧ)N�m��a��u��S��:�C�6�6D����*u��T�$��ي������6��m�Mq��ґ��6�P���n4�A�bE6��o4��h֭�y�,]I��T�1�9���\�U(����;-�ś@����AIrb�Vz,�[*�V�(�i�V�hzkE@U��[f3؂B����7y��W��(�:@�(x�j R�*`����C�lV�Me泭��^e��Ʌ^MA�<H��[p�v�cm���Q�\O��ڱ]��b���ax�1�;KW��Xz��=�����۶Si!ƹ���T�F&��뎶(�t���1��Q�t�l�F�,���S-�q����i�t��x����97&�4�+nWř��.gfE翟����1��D� b�Qz^z��T�5a�@w1
�Q[��� ��$���!*&���
�(��Cw��Ѕ�jeU�ܑ����ޡ�ء�&qY�ܙU5!^W�C{�r�"�&��2�h�۩\j��Vt�ĕ�eBc
6
b���Qi�x$��^�����Z��,H�m`E��,W���&Z�B쌹�SHx������]��@OCz�+-&���"���I�	9�sl�v�&�W�C{�������$�V�x$�V� �X�n��+tXp)��6Ȅ��mԳ�K���8�k3 �/ � ��9T��~�qi2�E��9	9&��\��S,�IySb9�V��n���eN"#�x��Y�wq���2TԢ�*���=�Sh �uK�XB-�X� ��L�Iʇ�.u���Cl u�z]/���>���k�n'tX�2��f���Ѯ�C��UBM@���q#i�l��D7���+u|�~�JJ�5T��������w��hE�'�=�S"@O�
>�;��vS��/���9	9U]�׳^�8��m$�JI����Qy��t�����_��v�V��!^W���� ?~�NEO�ؖ�T�ET��� � ��mC�����w�E�K ��{ʦD$���\���k
�Wg!' $��祓׍MY9Sb܀�Pr*����(՚�=��c~���s���*�����Ur�5U�q-�]8"��9kX���۲ѓ;�c�[��r��9�a��t������|ɜ��_6#�ym��\v�i�v6����;[.�y�����Yjm�m%���Ps��}��݊!���Y�wy�{�����$F
�!!����*@d�{{�����~O����jU��t�zݦ�(��,���ob�%I�\u���| ��w�dar�J���! G� �P��o��hQ�F�SV9��/�;��P��=2�3*�S"�@ @�}@7�>�����O�M$J�ި� |@��*ϼ���׵� �d�Ԅ�IlxXp�׆1�Z]��O�|�B-�X� ��L�Iʇ��\����ѿ<�!ڀ]���  {Py�{��������Ff�{�w1� x������2�$j�XoPΡR*��|M�16
��	>UB��Y�!f��{�u_Uc��h��֚��* �'t����l��h�eNn(�F��*�$��:ڊ�A�A�T������UJBS5q�Ӏ@1>1���j��9��N*�H#J��31w F� uU`�ȫ���:���v�W�T ��@Shz ���1/#4�*V8ڈ���;8��sȓ��Q���ճr$�[���1�֌��.�f�v�6�E,�H�� $���z{��*HҥcwP`"3�B�H��y	���4
��	"yUPr*���vS��/�Uo��9R
ꄈD	1Y߈��U��=�__�Jm�/+�*�[܀��r,^�`Ѓ�
��Q)R�)bE:C�yU-����t�)�I�y4�n�3��ȶ�y8�>W!MQJ�oSs |�T}�!�؆�~�伌�T�]�����7�o�'�iIT�̀*NBw�0�EY��&�i[e��  >�ܡϾQ��B��?TJ*R"B��vZ���hFC�3��cd�5�Gh�*d��5���[��׉3Ql�5�UTze�I̘����z<8�d��Y�Iٺ�-��O8��3�,n���QQ�v0���K��Ѻp�`;cLX�v�V��;����m�Zm�r�V=�m9�^��B���I���>A�*��I�g�qe;iZx="� � |���j︃���L��!#%�}9�U���2yV�b#ɖ�E�`C���u
mC|C{=ZN+����p7qG�=����87�Y3T���:���%���p]sL�4�8ar��.#4�U.�����>C}B��.��H��7�@�;舁��o�V��@#�e�RJ�4j�6��B�Q���L��ڪD���" ��0��C��}�/ﲀ�=�P�*�$S��!' $���<�6M�����7+ϊ^f����ܜ�2��M�-�L��"J�C~C��߼��V}�L��-`� ;���T�(DC�����r�T�X�
�B�
�� ZmIU�$$BF2BRJd( B$H���`=�"Y"�!P�#`�Q�@J<��X�e Hh"�G��LM�7 �]�Ȱ�B윙�5�4�'!Ѥu3U�EhtE��"�J�9G\��ucQ$%%C�z�w���vww6�� ���fP�&�A�D�,F M���؞!�R��v��P T��	�@M��%��I��zE[�Cw#�w�u��.��H��7�>����y���;�p:�*82GC�%�\n'Gib��zx��MR��$h�p6�x�6��7�;͙8SmT^� ���!�$�g�qe;i��C��Pd��|hm�reTԉ/4��ݜ�5�
�z�[U�S;ؽ�S�SIIX��� �!m����9��<	��TH�ژ�4�#j��:��&���9.7������n��= A�*���96������f�sڜ �{o�m
����RU#3q��;���ƅ������T��Uc������B��G�u_�OT�U�j���DE�� � *@��;��3XW9t2UU]ok�U���]-.���0�!�.�8��,T^[tfú��5���9wv�gBm�ڎ�Ʒk�,����ۃ��d���n!�K�$S/��i�&�iQN��yX��b���;[1A������w��F�� �z�6�n�4\[��g�5n����{�����
2��F��kQ���8F�P����UJD�W�/� 缀|hSj���H�O�M$%a����ڍޡ���+����`ou
�(�� ��},zW�T�TՎ6�3�n�oP��H�7��UF"G���f�Q�(H�nQ��cC�)�b_]g}u����؈�����=�~וw�R�}�X>��� ����j;�C��'�]U�j����A������ޖ�Ti#Uc:�G��wq@��=gA�L��"J���"X�3�@>4|� ��%I�M���8���%ٸ�Ԏ�M�vxcU$�T��� ;x�ާCx�[ �a��?o� �UI�I�	냊�k.�+4w�-�\���F# ��
��V.�
����#�g��vЦ�U���JT��UcwT�B�Tn�� s���LʢB�7j^ш�;n�Yϥ��T������"F�Ԓ��5U�~u7Ǐ��BNU׾�� �m+o�F�v�' 6�@����L��"J����(��л�	���2�$�T���@��9�)��������0 /	劇����	��<�&��'��.�%ހ�� ^z��A�@K�D�L��L�PR3u��Nx���������@�B���)*���mFgPo� �!�|,bjeH��7� ~ 缀|hSk`|g%L�IP��o��m��!�ٓ�.��Q5p>0O���P�Po�t�e;i[x="�ݬI�g!�V�}|в�B�$�Gm���Y$�	�iGfv�blF-�-�)H�t�������;U��Y9�c���7tlq.w���1t�bh똜O\h��ZŰ����6`��N1�N�Cn���n0�lr�v�4����
\��;�l3�MȘ&!B(���'1=ʪ0�f��eU)Ur��s������2�$�M,D�k"����d�|��S	X�B��| �@}�>�P���ERUSV4w�=�A�@;hP��FPT�����@"	sޠڊ�.fffh
��`�DoK��}u�G4��e�ݻv�e&�m<Dg �U&ٽwEN]y����A�<���!6�+� �`v �j=�A�@r���FUH�X��ί�o�:_Z���JUS"J� O�%������
����ܑJ�$%�H������'�.�Q�Z�Ѵ�ݵ����Tz�[l��݂oX�xB)���lA�*���@p>�t�������J�j�>�FgP��ޯ��1�#(*Ff�C�8c�B" ��0�Z"1h5Hz�0ŠLb�%L,��A�޽��آ�=�d�4U
Uc�:c/���B�ٜ��3	mkQ�Y�{�"�1�v�>����p��1����֚"Cb*�NX����i�T�Q����n"j��<s�ܯyt��N�gA�L���J���& ������0�A�D"�@Q ���H*�H*J��|����|���s�K�E0�6 ��I�b�(uP��P�!!� �@�H" " �۠3:N��U%U5c��fu#w�Uz�Y�k� ���cR1&ގlǗ1�US�ŋQeՓ���}}��	� �U��.)i����Yנ
	H*�@���!m�o�V���uT
����}�>� Ao��/zZeQ��U���`� � 0"�߾���� ��'�);d]��I�܀�r*�v���UX,�Bdc���$��CA ��	'�
%(�<Z�`��|)�4��#"$q��C�����l� �@ph�		�$��!$�AeD���1R-��`��ge��Z˪8�P��?-ޝ���vӻI0�z�v�<�4��ӳ�i�L&�fk���*�m�  8 @
P`8������ [@ I��m��     {s;h^�l֑p�s�Y�[kjVLg`��n�l�#m�s�n��6ZWf�]c�ݺYm�3T]$n�V�0H�cF��u����a¸Q������-p�aڧ��ם�c�9g�.&"q��ܠИQ r���C^�eI�qQ��٣V���I�L�<ۍe69�[!ݱ�V�[s[v+gV���۔Y�{v9d62<	!��ն����헆�ΪU]���n8F�be���D�������Fpٜm�s����\$�\tj���X��k8vq�s�#1�HR���*�5�-�8sd��J̚;�h���y�L��Ce)eV4�u�g�S`�v�rڀ�T�[k�Z����Ҩޮ��%[W
���)�ѭu�-^� m;d��j���o	�iMkd��6]�=a��А�{Y:�A�9$I{bR����X���X�.�h�a�^�������9�Yis	�2�*�S).�l���{W1�)ǆcS��U=eVU�M�d�di���c��6�8ڵmUV�*� t�C	V�̡��M"����~�{��	����Eх*<T=+�z?�����Q6r�0UU[u�j�vj����ɐ��[v�fn�k���Z9�@�	ۮ� :�q���f٬�X�㵶��˝�t�*�[X^nݡn������&;:�4`��{NѤ�9x��;�7�m՜�Nv�q�FT@�)�S��1UU��5PQ��z��ִs�ZxU*�]���`^����H&�=�����@ " ,��w���r�	X�
�(���C� ����#T�)������#� ��y �Ы/�ԙAR$�~��܀�ܑײ�.)i��$@vrERj���=we۶Ri2��hS[c����Ҽ�ar��TlR���TMp�
�(o�����̕y2��ѿ^��q"��
��T�4u�vy�,9��ٞz�צUMH%U�z�s����ے)U$�j�	"s�쑏^D��d�|��S	X�A����&9���ɚ�h����,�^�	!'р�l�e�6�j�I��l���	9�N%{=��2��fn7|�9� ڋ��ˊE�`��H����`<@7DU]P�)��Pߐ�=R�W /�P�P� ~�drwB��5(UX�j:3P��"zq��l�YE�VS���旣=eb(�x�/�[d�Yi�I�w��	胜��Ӌ��$"�n���چ��9-�r�B�A+{�Wq �� ߐ�zљV)R�5c���u�P��� � *�MHfx��A5d�I�;�"G����m�{���hAkLR/!��5Gi���x��
Y���H�vrERj�Ѫ&طE�b��J��$�g�qe;e�zD����*랈9�7�e4ȻO*O���ޠ�m�_5�h��H*EXoP�B�U&�u��*��"�U_oK��[�bn�@�$��8Z�5Ut�M��5�;d&=GRx��Z��^3p-�8��=V�D���w١��uIѡNg`�Z�qs��J�6$��<��(X��g��ܘ��q����C��9������s[�cFzT��q�t�;�k^�
^"[�7\�:��7M�.��ށ�o��E:K � ��}�P��v+)pe����ojrd_�y�Ǐ�-�6r���P��n����Jh�Uq��2�"�5���clZkM�S�U&�]��^�r�EI�q:�Pp�
�4\[�!FsĚ�m���1�Po��[ڪNU2/������"�f�<���
�AC�E��B��P�조�]�ZCg���^qx�U�ɢ�� �d��(��e�o���9W!J�5H������@n�D݊�\i��	�+{UIʦD2n����:���]pSF�3���Z�����çWg�0}�����{UL�L���ظ�CL&��Wg!2*�S����F6š��T؇g!z2�$U�B�X�)E"��"P(�!$Y��!P�@:�$�T�U����|��Po�:��(o�t�4+xd�ԩM\n�����S"
du��G�7ğ����p]p�,En��7et�ܤ5"��7N&�����y���z{ DD�!�KdU�R�ʥ��Hf���L��v+%q��e�����U=K�,_�u��&f�w�;�Q��5�����i��>Œ��TU�ƣ3�n���N�X�ֶ*��r���F����J[>�E��8�6Ц�UU�n�7�3��� 7����d#��e�N��7��S"�<��l����"�yRr��*��OEY�N!��A5k*tU��'��Ry�%��"�Zj��;ܪO*���zu��l�Ұ�H��l0<H�Skn Vk."��Wp(VL���s�q�F��ma:�m	��O.��^k<5���nN���k��ػ��>S�m)�bĚ6�n�%��Xݺ[e�!���qDk�����\eR���=I�\����������l���ē�����~~��{r��t��e�ydjH�_o��Ok�y��n1h&���' 7ܮĞBz/�/N5�JE*
�������F��;8�m�Yx�I�w�T�T��T���M�J	��oyT�U'�����&�	5��f��m�r<�dv�Ԅ#��D��qQ�.��q��N��Vgӈi��MZʝ�T���L�7x� KdQj��Pߐ�Q���OD2樭%�m��:*����Dn��'�h)37��;��P|�ǵ���J#IBq,(9I�T�R5c�[4sOc���e����N�����U'��ײ���ae�U' #���Q����H�"��R��J��<�w]j='^���e1���[R�B�_)�R��}��A�B���݇2t
B(F��t�B`7ga 	nZi$��#":7�"X�H11�@$"h������^�DqN�%a��H,`���6Pp�B�B7	RXaD"`��e�$))��3l���!*��������D�6�v�"�W�����P(j MhpU�K� �`�m؋��	�� N����W��ٶt�)�E�򾜫}ʤ򪞊�>�CM��j�T詍��@I�?P�������,"Ť�&�4����\�uF1�u�$L�ڲ�uW*�7�g1C�(�j��b��i6�	�P���O!�x�Z	�d��"U��Ry=g׳�D��M�N������wPhI���e �Xm =�����ƣC�8fN)RJ�!v�n��j��x�c���5a'v0�v�h��x'E[�U=I�=�2{���jj�w �7�����i��MZʝoy	�O!���MT��{�I�Bz*��ZK��-��:*���O*���ۣB��3��^�kn��vZ ȓ���@j��7��5���0U�,^�gmڨqü���]5Q�8�Է�.q�\ ��Q�t��9�6ة&m����FѸ�qb�X;���r�o��_\�S�*�u[Cp��\���s�Dk�Iʪ*��S�@�`��q�IL�wGnmG�PT$d)�JL�Ǟ��1C�!��(�Ô�0�ʝwy	�O.�߸��)��īӐ�r�yT�@?�#x��%�N����z*��}6����-��'!�
;��ƣ{�J�$੤�S5F���չ�*�Hnv,�n�(�U!(*E\nj���jbE�6�����7Ur���6 A1 5U��1S�Cni�&�V��ZM��lP{�� D Yy0�P�l�]��&f���C��ԞBdT����$4�o��]�BdU'��7���˷l�K-�m��P�{b���S����SU)
��&�9��on��2�b�9�UU3(*��� g��/&��1_L�zR�RM\7�0�d@Ȉ Q0.�L��s�}B���^ܑ�T���a�3SS�Z����GgY�DڥsR8[HWqF�ӹ0� �nId�R4UF����V��-�GcW*�����l)W&��R���w8�/%�7�,>��PT�"��:s$�![��̢CL&�K����9I�؏2�l+Æ��r�<�W��Dk>���h���oy	s�I�/�y���1u��l<���Kў�N��x�����q��[Gl�zNC��Ԟ�"��|Gʹ�լ\�����T�C���.��8���I�=�Ry	s�M�+��[k�oy	s��[�K�(*T�W���1��н�;Ͻߞ�~ώQ6W�;AUV���{U+�*�س�;>��ۍ�+�	Ŷ�Ja��٣]{5��gr�6A��-U\ݖK�p(GI��$�ۯ'/P\��lG;��{"��q��Y�-{.��m='�u�M�^@�wDu������m��t�BD�"��qrj�-�����/X6Sea7�.q�� �T(I�؏2�l+Æ��r�<��Ɵ��[m�x="��/�Y�Ry	=�Y�d]���NC��ԞUT�>�G6�)5k���}�9ʤ��B�vJ�[�Xuk[�ۮy�Y�,i+�-��e�;XY�9��O!.q��`��&�m`�� 4�� X��I	C�M�j�H�٩���ͣlO\�h&�V�����Ry}y���G�0��.C]�^��UT��݈�-¼8jNA�*��K�ksv�B�6N���m�Z�X��iG- �A�j�!2�d���ʷ����X�#���)�E�yRrw��jMB����~��A%RU�[��qX����k��C�?	w�E5����{�;��s�L<�`��T�*V8ڈ�y	s�I�<&���H�3b�b�M6p�ϧ&�46շK������i�k*NCo��'�9?�g[VCL&�K��w�r*��9�e��W�n����0}B\�LM�r;�UT�PY���[ηo�� �X�磘b.��!>��,d]��?r��=u'��?�~M��P��SN��]V��<Wi�>[���Qec?w��5���'����]�¬��RryT�B\�St�ipM&���oy	s�I�����M4�e	9��Ry�T �n����dR���2�@����w�_|�֕h�;�!"�d ��,, 1dH����kQZ�i�@<%&(�"H�F$
(@��P�P�B@��˱bXE�0� �i�F	�� �@�1�BF� J):1#!0
bIIQ�[���׮����O����n��pqv)V��<Ѹj�fpti՜I�@m[m�   �0 8���d� �  m� ��     �<�7-�'Q.B�0�[]qV�v�e���� u�����ԑ\�g(�d5�֖`u����v�@LXݖ�^UM�X���b�g��	YYj��ׇ�3�n�kn�Ԥ]r\�)U�8�Vl=t&�-�_�v�|�ŷE@�����d�OI��7s����ۃ�@\����{m��p��{-��U��:�W�
ݫ��u�0�5ڂ�q<��y7����i	�8 �)bv���Om���KUv	f�t��lk���F����LҶ�/�r�xnvp��t��R��lUGd^�f�ȝ�n������Z6�8/HM\p�n�t�JD������\d�8T'��oWJX4te�l��BM*��qΚL�<b�,�Us�5�O��j��� ��i���RX��m�P���8ٮ���,�n�vR���!��p�nrݻb	]��V竖�녮:�8���U�KHgGJ��������9H炙�j����`6�l�v�n�N��  O@�A�<X��;'n��ܓ$i ����F�iQ�&�ڌ���Wn�翰�0bb��'���	B�KP8!�.�9�&w/�J���*fgK����hd��8Z�aU�<���K��8m��5l:&]��G��[N��ړa���Hnw>�͸ 8�#\�{�Xz��ks�sv��!���B��V�m�xXcɉ������mœG�����h\������X���Uj (�DQQpaEH{up�=r�+���m�(�N��M�ܫ��%�4�/x��%�zD+{�K�jO-����g�d]��7�u��r*���92�ͬ�5��9�D��~�e7����@+3����}�$����EP�!I������|O̓6�n'Z^�BhT%U5���w:�/'� K�(*T�W�DyNzc{��z��@�~�S"�Ua�f2�
mF�P��ʤ�v��.��P}ʤ�.E�O��-��A��V��!멑&��L)XL�;�Oi��4Y�z#Y�VS�m����d]��'�w����x}-�&]����C����BdU&�� �ΆO��UF�ߐ��F`$^$JX��R��J�F�����3��{�+ª��E��}�V����ԞT����i���� �Dg��yB���phD�33@)��%+���y�d�Ȳ�t�;i��0��!���L���z#ɤ�w�u'!�ʤ��F�m�J	��oy	�I�$�OZm�h��9�Ry	�� ��*�`TC�TN�Ξ�99:���i�X$?]oy	�T�C����2]�a&����#�^��۪�;i���w�
���wRr��O.E�S�`%q��m`�oy	�I���)*� ���!ܞ���P|j+Os(��	������ȪO �<�@�wy�Rr���<���Z(WX>�n�0���h�<�����3t�	/5�؍P����"��f5C�u���뇶���;u�=�[%:�g�����b��K��3`�]њ�����݁��2D�H;'k�t��4U^8��b���IB��Ə��]�}�|��zgC����B:�Ӭ:�k*p�u�g���U)��Q����q A�������T��x� }���mi%�U.�L��!��{�L�����|�)�tcw��ݔma�ܖ&W�Қ�Sa��q @����|C����,��2��Ƭ��2��ۛ1����I2�j�YmM4ʓ��;u'�"����Q!�x2E��UP�X �� ��	�U'�z#ɤ�0�9� ���s�+C�ܚ��2�����$;u'��=7֛dZ/*NC�|���ۯg�����E�)$�I�"�x��9+���ě7��f;)3k���!2*��g��e0��I�nr�<��n���J�m��7�u�hM��@�8� ]�
���;�Ӧ4m4�K*NC��ԞBdT����$4�o���P��u�ߖ=�:�V*��ހ��E"b$q�H��'#[���s:���iK�&�~��*���Hv��!Ŷ�('�lU��BC�Rjg�G�M�.�ʓ��=u'�r-���}&Ք���myu�3�,��6@���W+ά몃��xU���u'!��T�B\�^��B����4jK�i�]��)�t`Z$��.4�W���wy	s�I�C�4m4ҵ�''}}Ƥ��O��̢Zj��5���mɨflG�H�XÆ���<�����o�D��H�_!.q�<��Wn��9���<�UTQm��U٪�[X��!�[k��E��ݜ[a��6����s��Z�/���y��n�N��4=��`:�aL��JE�u��[��T���'M�\���v�lR�ѝ����s�lmmh��G�=��w^�w|��]1&.�9����)z3�	�!�,���aBm�v��ϐ��5��EL}/x�ݔ���\�����T�_��i�3��2�]��~B��p��4�;�Ή��R���zE[�B\�Ry��M�ʓ���5'�r*헷w��h0�I3m�7K����pTlfa�W�he6Q-5vߪC[���W�y��]^]�Ua��>y�ҏf�Dh*FPׅ�{�S܄������$�-��ʷ���Ƥ�g�G�M�.���T[�}���6����%UQ��IV4���AȪO!���W.�v�d[f��Ś��[=y�����.29�^<*�c1���{��$�%ύo�nW;6�X="��!.q�<��7�h�w+*�O��Χ]Q��bP)�A��DЋjAM&�"R�N��8�!N���j�7���RĊ�,�5�$I+&q���eF͉0�� B,E�I�a ��{��F�i���}o��/�6�0M*'�pN�N��D���^�	қ�F�U@U�����׽̢Zj��5�������x��%�8jNA�*�N�j�<Tκ����2'�J	ۮwW��ݠy��=[�v��m�J�="��!�eԞC���	�wv�T����ԞC�*c駭6�ͬ�{�+��=��
���˯�V�Y���Y����T` �5��;A	�2>rw8U_Y*fe��j�8�l�� �>�KP�Р��n�R�X��M$�U����EQ�WSt��Fjev8��2p�|q4:���ƪJ���Uc��C��=�N7�.}4���Q�a�!����6t�x���D�-��-Ww��2�d�'n�x�ݻ�O*NC�z�O!�*  s���m�]17e�pry-T���ܽ�3uf�6��͜�K,�W5#�K�:�嗚�(p�m{k��e�����m����n����C�./i�`K��Ts�g���쀒�����>�AϘ÷����h�KX랚$��o-�k����f�7���c�p���X[��6u��="�<�C��eYL�eԜ�;�7x��:X!�K+¥*�V7Z��/ ��0�P��멒�����k�OI�&�v�ؙ�Y-��a�]�BlUw�YΕ]�(�DQPx��Xl]\�>��Z�8�iI����1��gq
;��8嘽r=骪S3d���~ ��"P4PC�؈��@�ޡ}����aNHUF�����C4��'�􊘓OZm�I��t2�{�zERydP��YL�eԜ���I�=���wj�2S���i�
_�{�N~ٜ�'�2t*����j38���B��ݩ���J�NC�z�O!�9�3h�[/C.��}��ߝТJ `�9����XN��qRSS5Fэ�C��7x��֙��#��f��w�ʻ����Ry�oI0�.n#v5�萫�<�e{t�Y�mZ��aBm�v�T����ԞC�*bM=i�e&��ª�wڇ[P�� @��r��U&��yt9ܫ��C�e�݊�\I��t��������_Q�d !��g�]��[���C���=UOqָ�b�N�v�iH�N��bR��rD�]mz�Q
U'�!���e�f9ͽP\WbO!�lG�H�[�WRr�U'��2��GqI�ex:E]�C�˩<�ӵ,(�U ��@�-9�@;�mE�=m�i&
��!v7���ENyB���|~m>Jda,��� $qP����L�ln����\���&ZEݸݺԜKѝWm��Zݬ�tz����z��ƞ���d�nڹ�zAR�{I�4n�4��\�%�ܨ��Rw�5� Q����b��͹�����m~��w����ﯝ���X�ܭx�֎xiym��v���6J�"��V���7�O�T�BC�Sv+%pe&Z��wy	s�}<�}��ɵHҕ7���}B�QO�֪J������ r��{�Sj���SH��8jNC���MCnq�I�Փ|�!&�L���8�WVzwC�kZQ	�An퐙I�e]��V���8�'��{R�i�v�W��C�
�Z8@W`@�4��;~B����'UQIT�cnC]�AȪO!�|�I��G�*��ߐ�yC|A���u���*��suC��W�uc���uZ�h<	�:r� �.L��q�{Lc�����ɴմQʓ���5'�r*i��(�]��\��oy"O!��ɤY,ej�<���5��IH% #dw�  <PM��[���Rw9�]�*���H��K�jO!�MI��B�9��Ry"��w4l�-�*۲M@�ޛŝN:�L���#�t�.�a�Y��!��� �U'��E�U�)P�S��o�P�R,����%pe&Ҽ�V���8ԞC>��d�H�J�@-�x�7�q`A�C����a*�*p������%K��iݘ`g�B�P�ޞt�,ѪJ���;6��<^�s������ʴ��l��6�c��}ʤ���'OrU*2���N ���L7�� �C����)*BMU��C�2@�����>����H��͹r��� �Ϫ:x����]���1ݸ}�,����~?�>����>Đ!��$�$�I$���@K%����_�6����T�+���g,��ow5��+���!畻j��%ټ�\d[��Q$DHAP�IEQِ�U�� ��"H�� H(�"�����Y���U(�Ȳ�Q�R$h��Q$OQA�k\��. ,�
��h�(�y@��QU@	�`j �AA
�!�B�UK�+�
*�SPA\��r*�AA�����",���(aG""�DV��E K"E AD�Q$DIIdT�S9՜�Jy���V�D�
 �t���:����{�I@Ƞ� 
2���B	��>�
�ڽ��W�����������=������Q����?�������W?�=�?���=�������z�B��)^���s����Y���s�?�����~����B=��?�(p�ڊ:��Y�??��~Oҟ����'�vY��5�{�>���������_�=��j��'��>v���u�������0���T�2)����}_���� "|�Ȫ��(BD�}����5�b}�����P����~�����Ҹ��?����|z�����{�x�H�J?��R�(	>(}?�x�hO��3��,��s��ϯ�90;���������nD�M�*��f�R0d诺�)��?��d�����7�#�N�
�5�5���iD����������4����$'���S�ơ�X�?��b"
�ת�'��C}�P'�
�
�9©	c�#D	 �FA	 �D$�BD! $BD$�HA@$B@!�@�	a �BD!d�B1BB$B B �#� ��,@�E! � "��B
@����� �"�1���RE�AR @X� D"!�! �H	�@��X! AQ�PH��@�@R AED@�U �@�  �T D(D@H �E"H� H�"�B D"�!��"#DA� �T��B �� `, `, H� A�"�V(� ��m � �A���B(�E*���A����@��F# $�0(�"A#`	b1D#ac`E�b�F)b�"F
)b(�`�`F D���`�`1F`1@��X)` (��$P ��(�b��D �@�!$ DX�A+�@�@BA,P ��	�� @BP!$� DBP �@�D @�$ �"�!�D����@���H�bE�P#0	 UPT;�-����k~�]@胙F?�/�����z=�^�f%��C���~c��>i@( 'm> �%�P�	!%B��Ѵ�$�^߁��LM����>g�!l>���}>��ߧ���}K�3�	9�|�6�p���D�?��:���G��W���o�������$�PAI��1N=�����=�~U�X}��P|��_�u�|����;��>��z��m����x���oã�I���}l�?����������FHW�����:�|������\��}��� T��}�쌂!_H~o����Y?��w��_�w��~oO��g�=߂G��>�2B��NP��	�UE?��ϓ���?g�_������U��i`�=�M���O��a�h�ۀ� ��	�����!�HPY~��/�M��U���֏��!�~���)��_ZiC�s�(�z<C�$�!�C����ԑT��P{������5��&t�����/�����P�����B�%6e4�}>�u��_q��� �O���
8}ʨ�'��~��v���!��_��G���,�.�h��������/�|���P������՚! s�����~ﴬ�~����}��������� ��?A���ѝ���o������L�*������ߔ��}�Ma$�,aIB}����
�����`l��Y�^��W������:y��?�����~#���A�w���GHv �<@��_�Q���r��4Q�^!PJ.���>���Γ~�'������������+֐�_��2���p�����L���Y��~������U�w��-�BSAm����#�9�C�%��������=�r����z�}�! ��.B2w�O�w�h�1���������C�?G��Ϣ����#P@O��?7�}�f���>�R~_���,���a�}^�j� '�O�����mDل���<�N�y����ɰ?���I���~��~�`W��l����~�����?�rE8P�ÓS1