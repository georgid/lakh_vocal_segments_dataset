BZh91AY&SY�p� 
_�Px��g������`$ 
�@D�	$@�{E5?��M����#@z��4�L�IEH=@i�     ѓ �`A��2`�4d���`F�b0L�a�101��&"H�d�I��j4h  ڙ4�dI����"b���?��~�XD@��1�է�+�.d��$2� +�Pg�1�9�~�DjubT:�hwk�g���pǄ�� �ҜH��
beL�$u���>�B	�N83L*�7qjY�q��ܙaT˟�o��$�x�� y}���W���4	�;��»��!wd<�f[ʃ}XOW�)�E�Q:a햡� ���^R��(�����M���z��C�cI�:$��`<`k��_uk�h�p�P�G�Ƕ�y��=U���� %S�WҮ�1l���ub뭻`�e�q0�1,OE����"�FA=E�n3tq�u��yydV��׷��r]9E�AԈ�**Z��q<MD���������<��@D�s��#�b��;�ع�B�p欓2�*��(m�q�3�MH��|#3'�z�s:3�(����{a�m_9�wd;O�Z�C�4�bвK�R1=b�kF�P�\X	��'��L��E�(à���rD�p �Q���x��BI��Oz9í�*J�m�s^��^ޙ-�QF��g)�`K���k#�f��[��G�<dA"I�IA������������ ż�W���	�Ӳ ��KI� "�F�,����
��eZ��PI	��-)b	x���c��{�����#�ℜ�AY
��}�~�nhQ�UL+��v�1�We�~��h�M��ޞ`Ӵ���Amy�k�b�E<�c���T9[�Ѫ|���+g���v�� <i�!.�@3�Y�=O���p�3�,���-B/;�!��t�|�<cݶ�w)`qF�"�S㪍
Z��N���ʯn]��v`_����Y=�]�]-�4Ύ DĂ��'E(X�C ��L�a�/z�>e� �Jyu���A��A� �q��7q�v~��NY�y!�h)2o���1ݠ�Ӵ}f�Ԙ N�����F��qd�Ě���[5)�;Y�:�H�sv~a�εH�\�r��,�&񿘃o����B,�����#S(/��y�PD�A�"p�Hw������\�V�!��wh��q�]���]�(�ؔUQ��������;v4gc.ܓC�fV�4�hcxi8��M��A�1NOyt=��M�����Tx�;��l("js��q��7Pb��s�?���iA�j� �c��:A=Ē@^��A����ßFg���!�Za �a1������gY)9h�e˟m��V�1�c�kL�:�8��W	TJ�c]D���,��g��FfpA�0�TX0?�>*l��c�A�3�X�ms�ns00���A�d�Plp��o�D�r8e���~��pV^(�ܑN$j�!@