BZh91AY&SY?0]���߀pp���f� ����ag~  >�@6� @P  U@ D� �    
      é)Q"�E 
	P� @U
 �)��BA)H� B�@(�� �P �P( T��<   F�#ѥ   d
����f=+�N��F���@tpE�9��2d�=�K�.c��a�s��ס���Nψ{ d 
Z{�"��2i�@.3@S���9��r@�s۪� ���'`��G;�o=��p} ��<��b�T>�<��k���� zX���	�WG =������C�U���q�����  �i+r� x�s�wa�����ip�H7��; ���8	�0��"H�ý�da�W�����f���`r�`:�v70u!>� ���
6�^���d݃������x	< d42v�^�2��1��ӈ�
8Y�9�M��:8�!��`�duJ/x@[P(���>���hS�.�a�A�@A���@$����U0��Z�=$���y��; �����ш4�����ѐ=       �*��R�J� h    Ǫ�US F  FC  '�T�T�P h   � S�!%"T �     �D��4�zM#5L�`�A���L�IH!D����a4ɦ`�d�LΩv�w���z��:t��t�ӧ|�E���� ��
�/����W�(��d���0}X���ݲ����<�/g�����'!�9�C�g����������ou�W�ȏ{��e�?�tĿ@�2*�\XI�cu]BBDCԵA��5�>�oJ�߹���}��L����
�۞_�%�1ַ�a��&����jR�c�S�D�C���u���s��t��Uf:t#އ~��;���h��w;���s�o�|q�ԁ�J�r]�!��e�CC�`���
`��!�L��.8I�d*E��q��78�!���v��#���a�,ka��	p�ef�O����{��;�SlӚCֻ���&�w��!�曬]ng�{�v����>N\q��BFbd��UqQ���ܲ]�sg�N�p�2��9�F��$��bВY�U��)��)��.`�s~�7w�����i�̩�������s�5򹩲l�&ɲlG���p��!u�������C�i�?XtH=�ْh�����)��)���iwG����đ0Z!r��m~��N�5	���9�>��L�y� a��}���$>�+D��3�d�\�Z�H�q~A8_|s���=��C�0�&Sxv�a�����s&D)�0S�Վ����_�����N�-ϡ�̖��{�/M�[��5�����&���Lˑ�>��v;��H�����
0�Aɗ�J�=�}>M��N���󰟃�X󼽼w.|�e�v7���p�~��\�o�x�sZ}�R
�NS���sY�Ǡ���N�˻�to�{߹߉���s��yɹ��t����A#�w`�2�m.�N/��%���s����么�0>(7� ��|�C�w1���c���6M��my|��溮n�}�}��v�8�4�t�2n&l�}m�f ��1{�������-�!�}��|���v̢#�`�X9�2s�)����� ���z���� ����s��=M��Ú��[����7O|#��?��/A������2����g;�ē�����ztB��s+lh�aO��^aɼ���y�����Z=�G�o���)�!w�~8��yޥ�߿w�\�w�Q�f~���)���T�t.���������Qg���������&]`=�|wK�^��k��EA����ĝv�LA9��w7����8�)�S	L�k�*o�ywИ�Q��Q?<�0Ӭ��Ԋ��?v��{�v�ɗ"\��NfcS�%�gN�4���D����NL������y�n	�"P?l�����wxzt���;y���f���kg��1L"a��Ǐ�t���׿��M8�3�p�U�J�Ӛ�u��r����&ɺW��]����3���w2�N$s"Gv�Xﵹ�̣��/&�=�����X8$a����a�1ߣ酯�̦{����������!��D·Y�2B9�s&D¦N��5��ӝ�u���zw��?H������ Lq|w?gk�p�~?S���{���\�;��~��O�>��;��L��p'�f��r�3X���3�3��߷��!�'y}��d�OFk&�"W3���"d3D�1�$&�~����sNZ���>a�
v&��,�6��0jT��F\p��H��"d��Ӝ��#�� �Lppp�KpIF9P�D�`�����x��L�r\I��AΦB�FB���߽�{�J8ԕ&5 р@�?0N�aGI��������zt����%|���vs��D~�`�ݺ4��~3��˽��$d���i��;�^r����M�9�o�q�q��n	ۄ�.�C��;���7v~������ܝ������ja��LA$����$��b.
�����>��~|e�oߩ�6�,�6]s��!�
��������gٿ����^���7�.�;�3���sg����t���ᯎ�d�r:?s��h��v�8p5Ne7�߻<�q߸���}�������ǟ�{\ܾ=�ˣ���nn�^��#��gsO�[:@{��l4�����N�M�T;��>e����@A�H�ji�L\<�{B�NB�ɺ��i�x�愛)\��Vk�0s�qS=�vB!�қ��;K�)�;���?���S���^K���z��'��\��
�p$L6��ɲ�sNNd��0����>�:a�!�A�ϥ����LJ���3ާLO&�׿�QJ&DDٓ<�B`�8�mβ͑���v�7
�"!6�>�7y�w�6��=I�Q[&~I���M�UǢs�cL��<%�?����`k4���h�}��_�������d�&<=�k��M�.\A�>�\_׃�}�|��i�%�r�HC�ƈ�(����gCۄ0\<��H�ᨑ0ds�)���?o>��y��$A�c���C'r½�K������#���'t�8�Ws�wi�n��ޙϼj^�Ho�ܲ;���;8o7���owyx[y�����w������B�1"`�;�����|np��49i�¤9�/9f5���%�}�ω�븎��l͛�0���.l�����_����� ����{�:|q0`S6�(Gq��s���{w���뉲l8�M�'1Ź�
`�K�s���{��9Ӵ���rK���<8�K�=h����r��3�o�<Y!��|ъ�
k���Z��q�f��cl|���f��9��6k�7rՍ�u1�3�-�y8;�ѷ��kb3��5s�&3w��0S�W{o0�x[��;�oƾ�y���Sa*�;�|Z����<���{1��9�rM�R31>�0ׅ��2e���"��'9��hu;�ܗ����~}��$u/�9��{���1�� ��%�
���s ���d�.?e��8q͐��B��b�q��ie��Ď'(9Rfz㐷��8���E\����șZs�a�Y'w����%6�]c���`<w�e�ʖ=��K��1����^��b�lB%XB	,J)���%<�z�޷�9s[�C�eฝە����!.6�IG	�V���1�"
d�H�}~���]�Ō�s����d�I#�1Ȯ5������Ed���rH�<��ho-7�5��2��l���/�*u[���"�`q��_���'�����4��|�4+��r�����oN���{��}�r���|:�1�d��|w$�
�Ú`�4΍sVW�'N�4�˜Lj.(0���9`�⒃�Z\���*a�������w���4�!@�:S�
���A"�
�
������7�O���=�ܞ��3���eX@I"C�\�D�se&X8$p��9��A�����K���3���KÉ9�2�MK�fW
����삙!D���!fGds'��q�12a��2%�&k��;�C��{�R��{Jci\�*Gx����bD�D�L,�
`�qȈgƚ5�T�\�ȁ������D���\��/���z���?t�@$�j�B��Y+�Œ8)��+���K�%����u��W��recY�e�]���f�ܻ����]�q�dV$.�_�~Ζ�)g��9ݼcov���-�>��{�?���l�>�\"bB!q��G.	>
ԌS����ϵReo�*�9G�Sr��@���_�g?O~�~��l'S����t�L���'$p�"	�4=�����g�}�w���o-�}�iO�{�-=8哛�~u�2^�M���toy��ι��ԇfF�z��D�r	'%�������ܛ&��M�d�6L�)�뮓�����O�{�a\4�ˈ�jS��8f�7��N��CR�C �̎0���uΗ������o��?`^	���2x�9ޙ�ô��8���@`���rN�߃�����8<8�v�t����7�}w�9G}8�aݳd޹ơ\�fu!���r����~�ɷ��T��Kv�������؛���&��:�;M7�����8w���΋��y<���Q'6{�^r��a��r��dGa4L�c�18�b�׃t����ͷf�ɑ!�uἯ�<��}`�S��#0�xDe"q4CK�
%i��|}��0~#!�JN�6���u[����1t����~f���L*"�i�/s���~v��z��^�8[8�R��|q @��d��̈C#�ЈK�5��N��s���
h�0.�)�p�/=��s�t�K�ԃ�3�S���0��f:����S��.�x��KH�|�n��ۆ�B.�����PAPp\�#�:�����)�5!��@[P�r�f)�~=�� ��/W�?a0�B~�\sԖ`�xy�����No,�ɽ�M������!��?�<�Y"`�
a�3���;�����M{�<sy=�<9�sRf̪�3�|���M�d���_�u�Y�\�:����$�q��s䣜��"�l�*�Y��vw,� ��ekq�9n��y��Ad&k1qd蜰�1���0�4;�O?��3 ��ĉ�83�XeϤ@��h�9M�eÜ��3���E2`p��j�H�>���t{��l�wl�7Y�����S
��O��a\�H_C(l�A���Dޯr׹�e�G2�@ &H�\gS��O<J�YrXXu�k�4q�����p�'\�y�1� �&�k���rI��,�.8�I�Aᷜ7+��L���)~���;�������׍e��{�
�)�S�
`�~�|}��-��c5�A��L!���rf޵���D��͛�f<�84�N��^��9:qH#�ݽ��d��'G��vkF\K�����"`�0\����q�����h�ݙ�jך��y��N>���L�qԹ�s^�eL50S�ۿd��P">�Q�Hd��Ph�.O�N�u�/���}Cs��08���3.ۙKdJd�3�~r���y�8g�1ɜrb�	 ��2v���ĭ�������f�Hr}�766GW:3��U2L*�I���l�N�s�p�!@Ap@��w�t�S���#3�,��l���߭��_$p�߮}�����ҩ߯_s��~�9��A������Φ
	;
��6~�t�p�qLQ�L�MԘ^�I����9��s�L��}��~/����~9���d�SYX��  m�kh           �	 �$�֨�hh�˔6x�B����۹'m�U�Y�j���
�V����%'�����඀�nh���)=F�X=�CZN�K�2���]�Ƶ�b䁕j��X
�jXd�cl@  pְ@ �6���%����� ^v�Pn-��( Kn�9���1;�
�+[Q�� *�SOX�MS��S�1�4���g��%�	�7�l ��mRlڳl8���D�����z7Wn�Zݹە5:�u�av�õR�U�`�"���!���UK�p��\8lm�H�`  ��ʵț���_5��j�-�Cv�j��8���
嶽g���UeUj��RI/6�H۝�-Zu��墶��l�d�I@���VΊ�@�.�ֺ��ET�,��V�<�CT�+��]���$v^��8��旚�r�[��ڀr�d��73jX6��8�"�3�]e����ݮ�VV�ªմb.�.�m���Q ���A�2�+ J���rԤ��+���bH�h	�B��UEJ�h[���M:`rɡѳDUZ�V]�aL�����$MK���r����S�g�wVQ��8�q��p&9Y8�h	.�`���6Ѯ��ݕ����UUTp (	  ���    �m�  � (  m�`��@
P`8 p!  ��h h�[@  a -��q   	                @� ���[_       m      	�[d n����
ۅ#�ZqՍ]o!��;]Tm��+����uS�x��A�v[u�1�B�UT6�8e�E�(�@UR��mUUpF����η3�4��3col  w�i��gj��1��+ϕ'5l�J�������-����gv٪��*���23�{R9��v6��"艶*[�������  ��)#Zݭ`��$�TKq�7(Լ��W%f�ï)t��4Xةb�:�V��R�"�B��c�ي��E����6X���m�Ʀ� ���kv�nש�2a�1�_)�
�gY`M�s�؄�mў�]���R��ꕔ`�iZ7R��e��[7Z�_G p�	b^�Έ)8�`yr�K�"޶�:Cf�66[�Ŷ�8��=��\���8vѷ<v``(6���&�aj��6���p��4�]&iz��v�qu�S֒����0�*y�j#Mi���F���=l��KA�4�5��J	r�T&�[Z˵6� I%��Ӱq#���Ѵ�v��2f�YInv�:�l4� q0N��-�AJƣ�W'5���Ӏ1sR]:�   �  �@ p      /Z      lp 8     �A��m�     ����  �:�4n�36��m�d�9e��l�.���0,��r����c�h�����m�m�ml��|�F�0=ۥ��@v��
c�l���]#N,M[,mr��5R���m)�8��[GWd�K�����8
�ҹR(�H�d��ںm�m���y�[v�j�U]��v�: m��f�q':�ڊ	��U[m�ܪ�)%-t*n�0
��d�Q��ݹ�B�`�*YB�-#�5�8yT(8vZj�2v����6�۶6�/C UJ�mD��+̪��]��`AweX= 	����nr�*��Զ@I�]���_S�~Β�r��+����+[%�JcU(��A隰$[l16����nC��T�K�s��l�Fŭ��aź���m��G��J:�:�d�]�}t�� �[.��t]Hmsu�C�^ EUl�)	pb[l�!��sUmZU��ћ��5ٶ��$-��h6�2�wq	!��|�\$�Kns��f�6�i):N��̓%�H��U��f�R�����9&pa�R�jO�����U*�V��O=;��Gtk���CzfT7$����t��𡖵�5ڼ�Qm\�)�u���q��c��zH�;i�a�gMfk�3S�`´fk�c���v:�n� F��M�X.!t�K&ݛtKm�5uae��ö�(m��l��V�MR��RT1���� ^�+ �� ���IgIsm����>pp -��m�֓���I�0  ��H�����NIn�krf$!)zD�����n����X�S���.P�����U�.$��숳N^[�u��y}�L6�����\ޕeS�Rh�pn�.a��\L��@���� e��
�S���UR���-=r�U*��� �ք���ۗ�ԩ�\�E��z*��ob�bg�!۱@/6�����S0,hV4cM�UU	J�ݳ��UUT��Cm�t�hm�˩2�g���-��m�m��U,�ݵ����R���	]���0!��*僭nU�F�N��9"8�LF�b)�=Un�;;�>�A���ZRRi��`Z�����`	�w`  ��hs[�#m��U.��HH$�ev�ݹon� m���!	��n������m�#؛ETV�ig2pt�����5!�[,�]�evMTB�,����BiV��V������] L���s�5Z��n�*�jm۪��F��㧱�����l*�/-� ��޺M#�E��-J����U[�m��X�^�{bvd\�:rH�N��j�ڐm�-6�,��  �[@��m��  ��
����D��P�TY,���%� r����(�'Km�  �F٪��Ps���`H��4ڂN��mzn�k���])E�j8%���[U�k񱈰�m�b���0�V�ݣ֝l-��RGj[�tGd��M��Y��3U����m˖@��յ�;hx8�j�a�[����=@O+s��Xf�tpe�P���x��hI�dvw(����<�#V���N$���(�-��<���T�+useP��V�������n;uc�]p;a�0v�j���#)Nnvy�������>=��8�8VB��EAuk㏶��.�;��9�\u�U�*��lM� �   �C��klm�BUz�h�ib�e����W	�t�]��b�Yf �tT� 6��Zk��amhH�PsEJ������mm%�%������J��UPm�krp���VÁ ^��Um��Tsh�Z�g����U���M���i�m���9mU�pE��ٶV�wY�@����Ur�c�y���6쵎z�%������^�^�   ��z������  n�$ �ж� m�  M"dյ���l�$A�kni�m���Hm��.�̓���a��S����o����&�^U�[N1]X�v
�JKN��-�W[�ɂ�K�e���0z.W6�S��IնI��F�ŵ[UW/��mF�l��S���� �hoK�i�M��pY"�\���U�6�õT��j-��`�	F�U`�T�T�i'�k%.�akk�$��Xck56�Y@m�p�'iJù�&]�n�Z�7k����� ��m���� [%B�  �t�^�'a� �`   �@�6�� k-��Vu�xm�	[I � ��|>H 
�6�  M�n�S`6�fdm ���0  �  ����` 6�l��9W�C[p�m6b� l��6텵o��H �P� �A���g᪭���
��K���[M����}d���`  ��h6ؑC��v�Yd����qUS��`�s�Rq�В5�m�hk����v�ƅ�B�/^*ۮ�V��@^wۍ��@�d���h-�d�Hm� �H	%.8 ��:�M��/Z d� �> ݴ�޶�	em�  ְ   �J6[�@   �E� H� G$  �`�    2e7dڐ  -�� i���rۀ��8S��U�  ݶZ�K	0�[V�D�3a�m��Im�}��/�g��9���HE���l���մ
A��8�t�["rk�PP!��/l˳��K��j�v�^+n�5�l ڤ��   ��gG[mm�l�� �i6  m�n��ˣJK��lT�Sk��   �� c�H�B�L1��@��
�2��U].��� 	�m�  -�����&�fK/$6�$���Lu�����ii�T��� �'@@���`� �@ ���U�ꫨ
U����pH6���f�6�� �aqd��z�j6-���$u�B�ċh�лb'�tͻb�����s�_\�ŹAI*v�m���@ݶ�m��Ń�#NjgE'Nm�M�:�& � h���  m���H.Zm�ů�}��C���-�   ؕW�T�JʠJ�� m$��˭ր�6���U�U�[���}���,s\9z���[�>c $[m�m -� m$��m��  ޠ[@p �l��   $  �     8   -�[_��{���������w��
m��ey�Q�^'��sObVjԦ�a�^�-��bw�^B�%x�'|���s��d[��cb�K"9�&$n#���䃔W�$�Ktt(uT�.�N��G���-j�J�{K�#�iLk5hh�1���2ư��[2����WJ����l��=QxJ}U�Y�j/r�T_Qx��rIG�<K�$�ʏ��Z�V�[g0kl�����.���LXO��O�~'�͢�T�O��t�a�.��q+�s��f-qm��C�:Wj�����S��~�ʧ<��%j)�O$_	{U��1K��?*��]H�9#��D'��&�NO
f�JkI�Δ}���k��^B��o�̣5U��6��U��,�[6�C�u��EʋU�6��[*fܕ\�+G�'i�.����rmh�M�s��8�a����?P�Z��왦��4ZO�Tp��v�%_j�qV�u;��M�NTW��66�Z|�=�Ю�}��~;J�S��G����ď�P�ͻQ�>"�?"z��}���#�h��'�����e��&i�ʺR�G���Q~��?+ ���\�y#��}��ʊ�6	Ί�n��\�� 5g��������Ĝ���x��,*L���e��&ɲl�V&�52�%m6ųm�Uʃ���8�9�w�Ow������ϯ�@ ��$�@S�-�Msg��78�WK���Ih 4��Y4��S�\t�n�hY��Å9�2�k��-5U�e*v�w-���hN�vGҨW/,�q������,F����Y�
���Ȁ �$Cmk]���jY��7bڐ�M�D�b�8p����  ��m -�;'�F�/YtV^��Օ�8[��1n��:�l�UG�[�����r<۷7�5�䞽c`)��Q�7]e[Su]4d��Eݚ�h);.k�����7a�OFEBk��9�p��nN�P*ʵT���N���Y,�s�l�͝��p�`�;Q<���:��t���vSd.E�
d�{H�b*�uX����v��2�؜l&��^�_f��t����U�ٻl���p�p�/.�f��
�u�n�`�,�!'WW9�K¾�*�WY4\�H����T����{nId�q�gh�θ���"ni�=skN����n�/V�e�FǮ�2�s]��nQ�lF���nm�X��c�/@kq�:#�\[<<����ېlQƧcI�����mhh�Q��z`&��4�@�K��E�5�G1��e�;��c
�vs�ml9�qKg�����ݐ�-�����W�[t '0k�O%p�vy�dV��I:{���Y˝N�5`k;��k��nK�V$4�wF��9,i;���[d`%T'������31�Yһ��ٷ�бH���N�	-�zv'e�3u>���=��',�2�-c�SUR�M!q,36Q�*9��Z�U�D#�iXZW���1��L�ښp���Jy�sv��iã��n�컍��md�� �kw[��t��t^ҵs%.��y�-���y��둞&���-Qٳ[.��cH�J��ѹ�NR0螹A�2k12�p��T��4��{fn�6�zv���K����T�R����U�l!SI"�9f�6�yn�v�lR�<ڦ�wwce���00�a�s�fs1��+��DWث��JZO�S��O�	��{�W{����,2e ��m���a���bm�ci�\f�v�[WI��x��{-��7��g�S���;:�$H�ϝ�vG��e���Q[t)-��ۘ����6�.��:6��v��N]t��N�u�c s��Gq;�]��+�=��Fֻ�Ռ�О��i	����3P:���\ٞ�=UV�*Ȉ���ʃЬ�Z�׍�/`�Wb�����`0�w0�ޝ,��[ZQ�؋kjJ�il�+r�B�X�(�m��XZ�.$�nгss�k`|_d�>�����}��H���D�}[�u��3u=��z�$�DRM"I'�H��>̙��7q&��hf��"�iI8���D�N�ՙ3& ��'��w^�$���I�I$�"�igԾꉽ:�ǚ�c��E$�'�'�H�I�|��xƶ�<o[���5n�@#b)�p��;8��[t-̧^��ƹ3�1�ޭ�[X��Oq6��"I'�H�I�E$�>�d��y��=c1��_�B P� � QV��*�iI8���̛�Hf��ѻ�H�I�E$�H !m���ۤ|�/��li�,m��I4�$�DRM���"U3sj��4�S�M��H�I�E$�$�qI����㿣���y�)ʕ�V�r�.nt�8�Jݟ�;W��,k���V���u��!CF���Y���I�I$�"�iI8���̛�Hf��ѻ�H�I�E$�$�qI4��/��cN��ch,o��O�O߿~���	��>�~����I�}��nlZ�Ɩ�{����
���Um�$�qI4��D�3q�n�OX�h,��E$�$�qI4�$�þ�_����j�%��CK6U�vÉ;c��sh{n��%�c�ۢ�Sr&���v"�CO7F�"I'�H�I�E$�>H���M�:�ō���")&�$���I�I$�>��76-mcKu=��z�$�DRM4-��[t��D�7q<�Ğ���Y���I�I$�"�h��! ��  'w�}Y�n�A!�y�7u�I8���D�N")&���ǰ�f�k1�vM�.�8��m۰n�X%��t]�h��BQl����0.M&ٮ�\�1���|DRM"I'�i%m���L�ڵ�����i��$�qI4�$�DRM#���}���Ǚ�<h,��E$�$�qI4�$�G��f)������ѻ�H�I�E$�$�qI4��|��6t�6������E [m�"�n���������w���uXl�]��Ԅ��d�e�շ�R��B�Cձ�\ڶڶAVZG�b-e���Y��:[�CP,gB�v9��p�*�N��\���u��{S�AMah�zu���^&�&j݋���7@�Y����=��nW���aY�6B�M5ݐuu�L:����խ�|X��9gJ�ی�n^M�ũ�5��� �wtڷQۗ��Q�^�5�pi��d��{2���30�e�r���wl*�ͻf睪��'&^Ղ�ٛ�.�m=��Z�M	�ֹ�]���kk��&�פu��I4�$�DRM#���}ɘ�VcY�<�k�"�h�$����"�n�$�� b�1\��ho=��m�DRM"I'�H�ɹgN��ch,o��I�I$�"�iI8��}�͋[X�Oq6��"I'�H��N")&�������b��d��r��<�:��Es#��K+�cjt蛓�����Qt��;2%>��I$�I$��o�b�Z	b��,z7w�߿~����0�#j�3ds#m���Ye��nE77N��ԝ1�5^�i��(� 1�O�$�O���ț:u��Mf�$�I$�I$�̙�kx���{����m��m�I$����D�un��ƽi�nI$�I$�I>�w����%�j�^�3;I9$�$O����f��{;��N����x��h%�Cx����$�I$�I$��Gϻ�6t�6��rI$�I$�IA ��%�������i��$��r�&�LifC�'ym��_��ѹ������$�I$�I$���bȣA,ZŏF�$�I$�I$���v&�Owuhy��<]�Xcs<.�-*Q�
���Ib��I�萔�I�5�oӌ,X�k5�$�I$��A�oڇڮ��z���^<z�I$�I$����D���ō��7�ܒI$�I$�|���bA,ZŏF�M��m�I���?�$ f������4`��b��Y�|�I$�I$���-	�^=D���g�6"�s�u�vC��;��sy�����ík���RԞ�Ʊ�$���$�I$����5�71caki�nI$�I$�I>}��E� �-�ǣw\�O�~�$�I'�����l�11����k��m��l�J[m�W�r�m�n'��n7$�O�I$�I ��}��,Y�1�`��^��v�}q�6�G�k��[�e�;[Q)�n"B&xF�Dn�&5�S;�v��b�;h�yn ��!M:ZNhm]$���3K�n�n#<�OK�fnG��D[���c�U��;��4���ɚ(9ϱ�܆�yh��x���ܴ�X�t���zz7&ͮ&�v0Oa����u�YT������[Qk�7��ݝ���r��ݥ �f̦``wN���JU�"�k����4㲕�=l�H�6зN��l5���u�����v+X���$�I$�O��)��K�c���$���H�m��$��>���SB��X�k5�$�I'�$�}��)�[h=q=ǋq�	 �m��$�I'χ䉭ѹ�����XܒI$�}�I'}	,�&�evS=�2\�W�,��:l�hm�fؓ�-�ە��׍րR#�u�h�???$�I$�m� �s5]Ibc1ci��ӧN�7
��X��h'%�	ӧ�$�}��)�[h=F=׋q��$�I$�I'���"ktnfca=x�5�$�I$�I'�1L͋pbn�ř��I'��d�I>�>�4,ݘ�׭�Mk��qm��Y�u��mun�4F�����]���Y��J��ri�ɩ�K����\�I$�I$�}��)�u�B�Oq�׮I$�N�I$�O�2���[�	��o]��$�~�M�
=��`D�C�p��b�i�Ls0*���c8n�)�fe��ˋKun��v�^8���ǳ��m�ך���t>s{�U�����e��^W�]��4 �d�F����ipq�Ùm+�z��5>z�l��׻�Gg�6T��+��\�nng3Us�`9:n�c�"���gf04��]q�q4�<�c|7{+��sV�"H�\�&Y{	��࠸��M�r�FL�/�0�\o.��d�\�c���9L�Jjn��&����r6U��/�;ӌ����DDG����L\F�k[ޭ�.���>/o7Y��25����#�[]�Y���+�E��3���G�5Ϯt���~|�/�}��<+�]�:G���/�4+�G$W]��|���#�
�}$vR���|H9}��I�}�e��fո14�q�����<�#����}�{�I�o�@�� ������)^`��KS���o_ 	�����${�� 	���q$d� '�ئ��Z���ǲO��h�v]�\��4/b�=��6y
�����}׿��H9������=KRo������{��m� �x�$~�J?~���D�o�ɭз3	���_m������m�-��"Y��������x�75��xm�|����p>����1H�{�jc1=y�5�>{����{��m�������A�(�O"K���U�zd��k�������ݽ�oԵ&��o����Ѐ��>��#�����##���6<ט�m<�,�"�9�t<*���:��c-��q@^sK][��q�7����kt-ō����������m����� ADA�~�������o��bkqn<Y����m�A>%( =�{�G��{���ĐO�@ �$� �@� #�e�0{���bz�mÌխkZ�v�۷n*-c�%��@{����{��"�����jM��__��4YX��,�b��{����q�x�I@�I���>��y��qca=O^��m��� ��?�~��������E���iR$�d� �1��i��ۤ����'i7�#q$�n�V��N1��̜v��ʷUm�v�7���PAb�!��%�GM��O[�����[aƜ`*C7�����Ɛ�l�t�h�c�R=hMvY{]��y��-�b-��&��ߓ�6���zvA��Վn�#-iA����۞����I;,L�D�rkE�O0ŕ$v�F�t�m�W[!K���ikW�݅ݺ�vKf� �4��wlz5�[cf*�[<��dTS���ɜ8�u�5;ڎ����˸n~�	Ɯo�ض6lF��=����m�-�� [m�,#����bz�k�m���  @���p>���"�o ߫�w[Ʒ��3��m�����m�����|�@�S[�����O^��M��"�om��6�x�QV��cķ����-��> AD��@�����G�߿~�m��m�f�m�:3Ҙ�5���e��%J5�.k`́2m�k��,mf\�xg�&d�o6N��k��ݓe|��{�����m��B ~�~���j��n��n-Ox�k|E���<I#��A$q�Ą2`c�Y���4s�ƴ�R.��,S��Qi�����#�������  	�AD�����Mn�Ś���|�߿~�,���I>���'�����VeW^x���mÍjF���V*��k\f��k�����>���#�F{�3˷R��bz�3[�m���?��O�߿~�~���m����Atbl&�Տ1����[�\���t�ᢻ&�Z�ܬ���JWd�u��:fs��v�ףqkA<g5�#�����m�-��&�o���y��w33Cz��o�{��  ����{��m��"J�Z6�x���O_m�����}�  F�*k��}E�U����@��p?~�x��e�0^�KS��Ś��	%�"��߿q�{���o� {����ۭ��Z1����m�I��{��#�����m�'Фպ2�Ndd�n��Q�����vR�&�S&��wKAf���Z�0��s�׷a��Jm�������[-�m��[m�dU�hǁjY�����x��{��?��~���{��Ą@�W���{�3kō�����[-�E��"�od
���kq6^c;��#�/{����{����} ��@ '	ݷ��i�(i�ԳC��ko����m�����[m����~��Z�p�1�`�'�/=�{��pH\I�{�eR��P����?�'z���#��f�ŋ�#�����m�-��� � > =�{���W���ĳ����f���m��B$��Q }�{���{��?�������.�46��� #�~��f�Ѹ�/1��|G�߿~�m�z�h����1b11*ŭkZ�5����E�MWSOV�f��ź��QD@��{�G��{����~ ��@ �~���o�������Գu�ō��x �D{�������o�A D��~~��E������D�4ې�T�:n$WE�z$=U@l��[Z�SM�ŵ���}g.�C��f
Q���	��6���6!�cq�6󎛱��8��jv�m���9�l8z�Q��`�&v��g`���6�����km��Gn����g��lS�F�S���9]s�6�G��{��t�n���X��Y�a*+wX�:m��.��u��˸�au��n��\����~�3;Nr�[!�wwZ�ۖ�m�ގTӔ8X��ɳ�j��v�ܛ�A���ߝ�[��wbY�Fb�x�[�}���E���o�$�}�x/{��x7e�0�o�����m�-��6�x�򘲆������u��ol����@G����{���#����-�KR�׋1����������"�]@���{�Gڼ���ؖ`ј�^,{܈��ď{��y�{��-��{�������:ۄ����a��Ye8����=�C�L̛�6���<�{��Y�{Y��m��[k��m�E�����{��>�ƭ�I=In��ů{��x/�$����&ٴ��٫l�a�l�6ٛKD˚��f���UWr�W@�Q����������-���	ePyh�M!�7^,���{�ȋm�H� $@�=�y��{��>EV��\K0h�]�=�D�A! ���{���{�ȋm� >$�Q@$ @��{�ȉ��km��Z�y�6��-�� 'Ă  I(�����q�������|�E���4�OkIjո7w����<�u���Vz����X]�wD�l��58g��)�"�f�[��OR[���׽ȏ{��m��-��$� �������<�|14���Ř��-��? 
 ~(�߿~��~��������y��-���%�4f.׋�"=�{�E����JA `$A�?{���_��mY�7u��փ�a�� -��E��"�]@�=�{�G�SV�����Cm�o{��x���~���~D~����"�]D}�>�˙�-m����l�k�d@3 �>x�jָjk��'k����ou��6�g����Csu��m��������[k��m�GϡU�P��`ᘻ^'�܈����!=�y��{��-�� �mY�3u�ѭ񇭾"�]D[m�G⇽�?"=�{�G�[ZI�Kt6�&��G�C����{���"�o�pr�F R0 F�@!|����G�g����z�x���m�����{��#�����x��`�ki�Abz�=љ�f�Cm�����㇚��L�n�1��q�ݾ�����B��/嘳���{�ȏ{��m��-�� �ID{���#���g�7^��񇭾"�]@��$��{��=�y�m�� G恵��OR[���7�ȏ{��m��-����"C��Fn0�cǋ1��<A{���#����[k���^���#��^�Ř8f'���D[m�?Q#�_�~��"?~���m��0M�$b�?�X~� �QP��k�]��\�3!��� ���9�7��0�݃�"b"�ɕ^&&��ؼE��b(��P�pq�Mǃ�cL��i����:NT\@��8�TrM���q�����͆C�d�$E�ٿtx4�	�E2I���&�k��ӧ�0�at��D��f[(�&��Å�S�A����H�e �s��&fc}�ͱ���M@\V��4��{���DQ6�� �_�ٜL���@1�I$��,�F�$���H9����Q�b{Й�zw�<T��L�P���yss S)�����swֺ��<��a�:ȹ*PF'��`�@'�>KJ�	�A�p��X>�����(9��a`yO>JÊ��޸�f�խ?�󺻵�6h��$p\�<�-��� �9��p;�?�}9�n�.�݄��� -���kj���:m�g;(i%&9QJMtή��U˶О�[���x��Z�ʖ�g\ �\�%�#Ckh^���ȕ`PŘ�cu������3��s�e�SϞyή,�vw#Ϋd7CI�lC��$1ohv�Flb�]����-� +��� $�  p �  H��[%X�;��y�������K� �n���r�hxu��P�V(����뫣ycہ�u�6�ltQ��:9�wѹ�^�=n�urT�W�ѥ��rT�8�>��/�+sk�S���h�glY�C\�p0 � �mҭUq�;(;���nx�X�\77�lÒ�<j��j  �#z�,v[,v,A���J��r�9�85lgj��`$�����֯N�*']�Qp�ʪp)A�7\c��cn�fH�a����nm�H«Wrٗn�Fk1�0�Z�� 5%n;lU8݌ֹ��/-�\������n~ꋶ� ^]��wn�Z�8tv�C[q���$ֹd��4���Q�ƴ�d�"#�ۍ�ة�ٮi:��K�K��D�rʻ�m�m)��<nÞ(֤O�����ݷ�� �\����ۤ��{U9&�T���F,ݱ+&�E��,���k �n5���bs��k"	<�,��&��n��Drd�3$���۶�L�og�����4fI3�c5f3�ԫAm���a�)�i��AӐk���֍��չ%��^��w��vwX7M��0�݁�5t�vvUg�
� ƞ��a�5pb{Sj�VU�N�ݲ�$l��C t]cn�u�ƻi:�;H�Z�J,Ì͍>�+P��V�ہ���s[��S �i�rFq��C���nN�s�R<�ku�cj�6ĵn�g�^ʂE�pUt�j+o�>� ��c ;K';s6iYe�2��"+��X�N��0��.!�]s�]�kU�x�8���KU�<��-kJK����A�эDV�M�n����`�n�>y/�����S���ҧc����_�^��S�{\H��8����yw᫋���p�es���U�f���&$\�e,)z�	!�Ѧ[g�m9"����l�x�̼@��[�����l6�)��u���W�����Gf���M�1U�pݤ����+g��|5�,�k��j��ln�r�\t�OX���{&N�닙VZ��'[w�?o����Y�v��ζ�b˃�[r��%���L��\�D�uŀ�����Yy��w�v`g0�9�6���&�ݓR5�7"nx#b)�s�������c��bM�JXmd�vI�>�?�:��ffn�Z)�[�_߿?"-����$y�)�{��>����$�%�o{܈���� ! "� "B �~���D~����"�]DH~գh���x�f6��mum��'�	$B({���#����|�)���.��]�uמi�ՍS!�f�/{���z?"-���� A
%B$�$$@����G��,�fn�Z)�[|E���$�B@�@� HD�����{���"�o��W ��i^��.捖����Z9�Tdʹ�ga��w�uζ���)��ei�1F��Q$���������Cm�ǽȏ{��m��-���B�������o�n0�cǋ1��[k�x��?�0��*0˧V<Gu��y�y;�0�i��3�:뫧��kϞ%�N!�&51�5&�a����~���"�oĂ��H�� B P�%=�Y�3`ᘞ�y�܈�����E���#� �A� �D��{��'���G��Ve��z�6S���<�D A"}�y��{��-�� >%QD���qg�[�z�����{�m����Q�x�mu�I�����9\�p�65�<�]��ص�5՛p������۬(\��n �&9ڏx��]�<Ǐ�o������m����W�I ���D D߿~��O�=�Y�3��1=y�w�m���ED����#����[k���j̹��V��xƶ�m����?��/���x�B������CY[J�Sm�ڔY� ���|���~}�-�$���y�w��P#����߿q�~��"-��$x ����Dz���o�kКǏ�o��lD~ � ��+����G����"�o�>��n���kV7�tv�y����N��y6�����Q�ɼ�G@w>���٘�.9����o��x����m���D��IE"�����G���n��hl��km�[k>!��@ �A �G����y{��"�o �E��(����V�����o7��d{�������ĀC����y{��#�?j���f͎ۻ����O�0L�0 �	�
��~������߸�������qf���٬�O��'%?*���Yb���F�����>q>��s٘�㘞�����m���H�8�-d�T�)��L(��?~������߸����>Y���_�';r�Z�����'#RRqs�o=���4;��<Z*v��4�0��z+�}���m��m�EV��
$� A$���&`�A��f� =�{�G�ኬ�i=If���v�d[���FV4a���&l)"$AD 
>^������q[���[ed���6&ե�g����ס5�'����{̋m�EV�ȶ��|���b�K�bz�;����Q�+MC����?����~���m���% Q)	���y��yf{��Lhl��km�[k'�$Q���q^��ȶ��~A]�C�ہ ���S�Y�l,^zZ3��7'=[�P4F��,�7�aF�ݠ��nd�`�Ͷ6`��Sn�n7.��:.�'C�C�-9����	�̇OpݭҋrՅc&6��`	��F{=NF�g\����@�<�BvR��;����F��աtR��<�)�Y�7T��ۮ����:V9f��u6h-�i�q�[��Q}]���w{����5HE�M��<�$MǕ8�A֒R��E�-p/7n��9:Z	0��a��%���;_2=��U��-���  Q��@~_�~�ȿ���o�Z�&����[�*��|����{}�y{��"�o�R+�����bz�;��E��"�mg��C��߿q��߿2-�2�����m�#��z�̏{��U��<�@{������*����%�����#�oU��-��[m����������Ij�Vʮ���B#N���u;�*n��;
ilb�K�np��p�M��ůk<Ou�#�����x����-��jɊ�31q�O^gg>d[m�I P@��GNߌ�d�EV���I#�#���3��m�Z)��|G����̋m� _�@#�~���#��߿q���OR[��{�Ϙ���{����E��#�$"�^����B{qo�k��Ǐ�o���Y x}�{����"��þ�E��6l�$��JE�v]�F�̼6��\������.�6h����9���4�d��H����}�[m�m���xy H�{���yf{ۭ��M��m��o����߿~�������"�o�@�YC	�Kt=��7��m����YD�
u�Uf��!hg��쿡B��C��|�>���dX��f�Z����]�w�]���TY�%�3RX@_�g�ߴ�߿~��[��� �{��,X��س3���]���m�O�%  H
${}�i���"ܶ�����n�m[��vM�����nS�&�"�� �w����k�fP��8�8o:��ۻ�q6S�5�����?~��[m�-�n���{������Ԗh{��os"�o �"�	�{��#��߿p6�x~ ~!�C��-��S	<z�=��߿~��[m�m���x�* ��3���,��Ȅ���p>���"�o��/�kY�����p1�j��8k��me�J�-�ʜEڋb�j�[kZ��kWL㮶ۃ{��)��޾�om�����[o�������~��?h^��.��
���/=�ȃ�e�V��d��Ҳ�lhn]�3y�=gM	�Kt=����q���"�md[m��P�{��ꇮ��ũ��=x��|���{���{��-��� ��,����,���1=y�7���������"�om���\V��hl���z�����{����p6�x����߸�߿^Y�0���C�|��q[xm�E������<�%�]�h3#�mNU��.98��ٳ,0�K@�`�����mev��Gl���mh���?H���X���v�uYd���[b��Z�Q��ïb�K%�α�{n�'��.km��!���0�\f��np]:�B����^9��ƹ5/,����\��Ռ9�ͫs�g�4�Ga%��/�ݺ�0g�8�<,q%�!�cu�za���S"v�|j#��\n4�mR�v�㓶l6G<̄�޺o!�-�+ĺl������t���2v8W��������:���y�c.K�ʥ��Й����M�[��D�<O7_�3߿~�-��6�x�m�E�.(.nn�.9�5����-���  
�?�~������������?x~��3u���Z�6�߿~��[m�m���x�h���z��[����~$����߿p?�~������~$������{�{ږ���x�<�|��"�om�����|��f�e�m��cz7Nf��ڦ�)��ni��5���WwI!Ia�I,k�@�����;����\sk���_{��m���{��{��-Y���oV�V��^��o
6�f�Z�@n�P:�����\��6��'mr�ﾮN�Nβ��["yU�+�����8�[�[e�A����OR[��}��q�xm�|H!{���{��%B�Kn-L'���Ou���{���{��m���!{����ye�|�ww1q�[��s�"�o� ���q����o�옷nf��cCPz�`h&�лd���]m�Oa8��rMuv'Qnz�]ۜ��խ�����m������m� �x���Q]x�Ԗ�z�c��D���m�D���o*
\�6�x��-i=���m�-��F����@C0
Ɨ2g5����vͺ���v���������ɸ��s���O~qԾ_��N�]:�f����p�d������!o�H��,!\[�9��snr�cm�45��s��_NWɩ�����q%6��lm�߫��+�������k4��?N����۾���28a�hp��2�d�]=ds*�޼wٕۗ*�V�nG}#��mBc��p�&s<�LΩ��8ssV���9�|�(�N|�}z�]G<�q�g��m�gz㫷�J㮓�5�N�o=�[FM��7箎���w�����ꃵNhs��I֋uY���a�����S��S���`��^��)�
x���}��9bG�G;�����>��Z�d˙�����-��9��@^�������[m�A�{��������c[+F1���om�����[o���������d��6ɳ�E�E�";B��u��Hk˥s��id�&�ݕ�sS�;�`�#��^<�ԷC�����#�����m�-���K2V��kZⵦ;cX�6շ�ՋZOu�6�x�m���"�o�@ 
@Aye˞����\s�������p6�x�m���#䂬˙l���I��� X��&a��#�{��=�{������@�<0�t��M���ǚ��u��u�����B� �� ���q��1y{^<�ԷC��>�-�� �����G����{���m�G�H��[�ۯw�z�m6��h�n�v ݮ���**رc��Ld�sN�a�jSd���v��9����n�-i=�������"�om��-����2�n��.9�u���$���� �Q�������"�]D}�E�s7q�l����~ ��{�ȏ{���@H�>�{��=�{�E�F(��y��n������-���H���y@��������F,[��Ks5���n[t�m�E�m�-���IAHE� ( 	E�K$BJ�5���	��.�H;��&��:zg�n��`	�[m[d<p���h��n���mм.ŘM��wy�������7h�1�e":zsgR�ո�:�f���حO;]e���T�mnɺd<��Mv�1/�v95>LWf��!��q�V٦���1��VMFekm�����4?c\�Ɛ�'H�vܝI/���K�{�vK]�4�S]jջV]#7���@7b�)�.�-�^ݎ7ja�=��2���i��$p��v��Y�7p����mf�N�m�<�tyy�G����-�n�m���$ =����OxU����z�+=m�"ܶ�'�$�����{=�i�x��b��Ǚ���{�oov�m����E��Hnۇ��\%�jijŭ=���m�p�m�E�m�-�����Y�����-�ov�m��&ܶ��x�rۤ}�%�-c5�nun�o+�H��]�#��r`�ѴZ_3���:ph�t���y���kA`{���-�n�m���-�@�oe����n����ݤ[mბ �'B	Ďr��qX���� �?��>�on[t�A���y%��ՋZ{���{��-���H{��{H���q���Y�����-�wv�x �@���G�����$dI�M#�,�fn�ա����n[t�I}�{�G�����m�D�ܣt]{���׏.��d�ĺ�E�=]�A��t�
�ᴃ�����z��n����ݤ[m�-�nm��۶��Im�ՋZ{��ݷ���[��"�o �.)Vn��.9�u��ݤ[m�-�n��"@Đ	�HH����#��n���]ź�sCK=m� �n[t�m�E�m�-��m	Eu���Kt=�7��H����"A�{��=�{�E�m�|�G��s��cT:n9�<	��4u��C���q��(\��J55I3K4����훽�n[t�m�E�m�	�(@���q��]Y������3u���H���[��"�on[t�@ A OxU��[�w44�c���=�o��Km�%�nm��߿���Y�i�v��r�B�"E���#��~D[m�? ��Q%5h�%����j�NI0p"�9��I8H��o������nQ������-��H�D�{���{�ȋm�D��у5n\{��Y�y8ܻ:V�iN��G4�m��ͺcj�U�s�t�g������ٹ��q��z�{��x�mum�����?"'�*�n-׻�X1�m�ݷ���[k��m�?��{�-_��X��[x�����߸�nۄ[m�-�n~!n���L-�Z�<o�� D ? ?�~�߰�߿~��[v�"�o&d��\��ĸ�n�Yϰ�m�>!�����{��m�p� ?��q�����c�v܉�҆ܝpF�0�bt�u�8��5m:�1c�چz��x�<� ��%K�E�mm�&z��vT����z9(����"� ]m�q�bf3�Dd��,�]T���n���x��d�v89�'W���������m�u���>��6������z�qI��1Q=v�=a���&|�xr��@�K�6I)���mѻawV������v����ڬ;Zp�tqs�%2]��z����\���c�$YG��*m�#ޛ�a�x�nۀ�G��{���ҷ=�Ɩ�z��ϰ�m�?����"�om�p | �{J[ᩅ��ZǍ�����-��ݷ���I�&,W73q.9��Vs�$x�}�{�G�����m�� ��o��K�Vg�7^���Zz�m�p -��ݷ���O�{��)kLu[.x�8A�\����!��5wGWWv��B��F���O>� �$�Ų���ϰ�m�E�m�-��&۶���Kh���ŭf=|E�m�����C�!��41V����uD�?����������E�� ���������ĸ�n�Yϰ�{��m�p�������{��{����.f�պKCi��-�nm���%�H6�x�ﶕ�u�X��[[�ݤ[m�-�n�m���-�DO�в�ź�[A�ޭkt;g��e�CZ��e��u�3lvQ��t�]�s���sҷ8ja<ŭf=|E�m�-���H���[�f!�nf�\s7X]���m�? H����G��{���GϴU�s7^�яci��[v�"�o$�v�����8������9�i������?�i�'}���#�m��-+r�ı�����vm����E��"۶�b�[�ji5�Z�z��nۄyHA H���q����-��~�H)���4n1��Y㩂��L�:�ͦ�I�ͻV)%4�Dܶ�W7Ad��[�����39�m����E���(�%	�����x{3=���n�x�M�"۶��x�nۄ[m��
 ( ��x���X��[K{����qݷ���[v�#�BaY�m�w��w��������K�5�i�H������~����"۶� ��(��#h�R�[���?#?�{������f!�nf�\s7X���E�ׯ^+R4L�+�%��k[kXG�߿~�-�n�	k�-a����>2*uŐ���n�a�8N��yIl�z;y��f=�כ�ff6�|E�m�-��ݷ���[NL���n�����vz��׍��,�K+�ֲֶ��k\E�m�>�-ҷ(ׁ43Z�z��nۄ[m�� "E�C����G��{��2�C*���\s7X���E��"۶��xD$����>�fg�V�c���i��[v�#� �{��#����?��������G��ui�	��|�?�u��u��u+|����W��U�ʹ;77;�ܮ��C�$�י��9����f�f��Tr���q�n�8��:m���.���=]�7�^m����e�@ [l��.�:�/'Ok�*�n0q�Z�l����J�����u��6�̛�s"��p�-az����/�U�5���.��:yܨ��@#�|Oeݗ=p�=p�ÑU�[��zM�k�-��!�a�y�}j�:�r�֤$���6�!�u�q:�  ��  �����9�[=�U���nK5�4�m2;vT�XR�u��(��ȵ�����v�b����1��y4�9M6�d�/^0Ş�\�S�d��g<$���5�6sh˙ԗD M�ѹ9���4���� ��@I�l�i;�:D�r[u�X�����s�Dی�1�� 1\�eri	ں1+[�e]\�e`���j�hE�q�g&蹺6���M����s]��2��l����Vy.�
�J��A˶�ڃU�烄-��(�'� vŷ:Lv��̇\��"��6˽��n*���J��&Enwp�Ǝ���.�؅��ut����\��*�y��bꆂ�����X�����ܙE>ѷ&��k��c� ��HLVȸ7k�z�sTݽ��B�MȅD��WL��8�W ؍�uju��
�-�s�
̀�-���OH�N�2�]�.�;q��'a�e�̸wmqՃvɏ+Wf���ɳt�Us���MHP�O"�<�ULXT��^t^�@Wq��k�Z2J��m."Hn1ݖ����ٮ���[l ���մ:�,��2�`�r��l�W-�'e�.t���cZ��l�iN��v�6�\��I2�-�(Ui*'k��K�ˀ-�6��e��3�ԫ3�h,���e��ˑ�a���m�^H��:iѷnI��n��AT� l��d��ݷ]6 5�X�9�f�b�vδ@p�������6V�u\�N*��gus�h낫�5 N��P�d�(y%�jJ�����l�����q�y��Q�Z+�0�4b�svwl�ZM�l�.�ZK(�4�/&Tܑ�u��Gk0m��Z�w\�ͲK��l��| �|`gP>��e����UuI���@yTs�U�<�i_�?`�i'�륗[n��7,�&�1��J1�����#�dy��\ڶڶci�癁�����ۺs�t�-�;M��O[�⭝e��6�ɵ
�5c�u[�l��s�1<�5�z擧�\%Ɋ`������|��7T�h���6zF������y#��B�����7X��WKJ��R�������e� �m��e����h4�m��85X�ev9��̥�������F+t��S��:tZ�5�x��j3�)�i9��x_1fn������#��om�p�m���AA$�>����%{�熼	�Z�c��[v�"�om�p�m�?���I$��f~�!����b㙺�g>�?~���m�p�m�E�m�>}��e���cx�5����I�FP�	~��~�?~���m�p�m�E��˯f�[��iowa�x�nۄ[m�-�n�	k{�v���`E�����ώ]!�IN�u�c�&<�N|�]J59��f`����&���.�5�ZǍ��{}�"�om�p�m�E��bV��b㙺�g>�-���A?��v0j�a�\�k�\�7sL]�gZW���c�r�QL>��9�ժ֪�C]zl�G���"۶�e+�77��,�m��[v�"�oBP �D�����{��%�L���n��o�vm����E��"۶��A[�r�M&�kX�"۶�@�E@I{��������m���Gۡ`����^�5�a0%+����ӹg�lywC�:��p<� y̧u���1�*�����ǻ����[v�"�oyD�@�{}�"_
��F�X�K3[m�ݷ� G����{��{���[NL���n�����vm������"At�( P�塗2-�,�LB�L��W�s��/W���L����q'���'�����Mbֱ�|�B�����{��-�n��A ��{��W=�����Y��g>�-��]����[v�#�&J�.{^�cX1�UF��h�*�naq�B����CŐD�k��t�X5'�75�Y��o��{��a�x�n۟�D��@{������;��x�4�C���wa�x~$}�o��{����nۃď� !}��[����X��x������������{}�#����}�7j�3�V%��י���^���#����E��� RD � �ۿ��(�\ѹ�PƂ���|E�m�-��ݷ���~$�L���7�sX�n�e��8K�#��n�]�n���k-��-.�����Ms�=�n�;6,մ�u������߿qݷ���[v�"|(�d�A�Z�<o��� ������ �>����D_{��>}����4b\pfky�܈���[k��m����?"'�P^���,����?�^�������q��"�o>�VeǉcKt=י�܈���[k��m�E����t} @@�		�? �d2�+��	.�WuxCF�����]:j�f�I��煅�oN�5mD�ɍkk��Kn�,[�]��x�v�It��D�U�%E������km���g.8yT����-�2(�"Ƃ������G4��q��z^k��;u2��s���ۧ��kk(֩&
���7Q���\JY�Q��a�dM>�`�*��.�����)Z��.�kM�vt7���ܛ���iy�@�����pޮ���&H��NR}�z��9�����뭖�݆�:]ݭt���sI�Y)]SR]n���>���m����W�����}�v�`ǚpq��o7{��x~��}�"���e�p���.f��z��f�m�ݷ����(Yv�-���)L�K`�՘��B*�om�{���~$���o��}�<*����0�֚m�ݷ� (��{��#����E��"|���~�9'!�c����{5�۪\�d�I&�H�89uλu�zv�wl;8��}��|{�e�E�m�-��ݷ�D.f���,�����nۂ��G�!$�$x��H�{���G��o��m�E��Wı�ַZyϰ�m�E�m��@�����q����>�Ew'���f��o���E��"۶�Kx��&�Wvi��f����E��#��A�����#��߿qݷ�����Z��i��xό�^��)���9煪5�jy.��ܺ�6D#���Z3B�x��f��������E��"۶�Yx�e8����c[�'ϰ�m�<@��	@@~���a�~�����D�(�*�ǉ��f����[v�"�o��!��������" 4$b(�9�Er�	E�l�ܵ��fs���s��';?���R({~oϸG�[�"|��\ۨ`�7^,���$��z������e���/{��a}ꇳ4,׈=+7u�|E�m�?( P����G�����m�GϪg���O�F+t��4S7a3����ѧ�f�iX��)�k9��y[q���f�\����[v�"�o`� �����>,�3<10�֞���nۃ��@D#���߸�߿o��E��"�n�pc�C8��׋;����Yv�> �  ����#����G�"
慺��f��m�p�m�E�m�  � ��$�z�q-�1\31�ƛa�>�-����$a��o��G�߿~�/����{������F�3�8yx3��!Ë>8z8��%0޻T���e��\�GR��CH�d�GRhf����[v�"�/m�s� ����`�4����=x����m�<@?�# #����������G�v�#�sB�x�4n�m�ݷ���[v�"�om���Uf��6��}�x �(/{���{}�"�/m�p�������M&�kM���nۄ~$�F�߿~�?~���a�x�>K�u\x�jx޻���n�i���iE,7Q��i�v)f��[����$�@�9ƊwX��jk�S�ct	�mu��$�k���m��.ƛ�uE�\l���q�8�1�D�r�V��3��f:;
�$�r��.�6��ZIX$d]�M�؊�,A붰�̅��EY�=�m���Z�h���Q�vF�b� ;��%�)ݝ��Oa���wa��X����G};��ڞ���a��@��� 'r�.�(���s�i����;�������`{�;X�����-��ݷ���Y�a��,�XKYY���$�0~ �!}}�q�{�D�N"~�����9��m�>�-��d�D�N"L��}Y�,�54�����y E�nm���$�$�q~E�i\t�b������E$�$�qI4��ߟ��w���p�j�ݵZv��Ist.bNMGT���P���c.�a45O��oyԒQc	6���O_�}�"I'�H�I�O�StU��05��=�#��@�$ ?H�Uۤ[���"�i�}gԳ ��Úֶ��H�I�E$�$�g�}R�7t�ev�v>��?@!=�{�EV�"I'�H���@��m,����"�iI8���D�N#���߿���V�D㌜�pju,���&��f����k])�����Ms�m�Vrq���[罤[m�"�iI8���GW߸� ��Ú�ׯ��I�I$�"�o��x����7t�ev�v>��-��I4�	�-���<�AA��!W���ݴDQrf�`��c�م�q?p�鉐���7[Y1�+��fL�X��3'tG���qp@~^9��y@SEQvfNd"Z�$��B[�u5cC\�{����u�}9�&g�I��&�(�AC.�^��Ò�Au	���	��¥ȐH�9�p�و�r��	0\6k4qy�J�q�iۭw�-^ѯ���[F�hک�Wmۿ6�Ӻ=�wOc̚�֛4�c1��2b�"���W2�l	�N�B�k�j�2�dˎ\p���q��:8{���v��9�n�32��\�ke��kgMqls;�&9ۆ�cM�I$��NN3q��A..��q�+���\�L�L��P��,�����I��⻺s��7~C7ww�: ��p��t]�է]quV��S[�}&ϳ�y������3��Bp��i�����0K2J̬�7Zɪ��m.w3Pp{20QApPC�=a	$�����a��9����-�H������G`�ڨڤ�|����5S��4A�B��T~�˨��#(�?P��G�$�Ƃ�@�|���E_%�?��!��B�[K7u6����D�N")&�d�q��7�U�V��[罤[m�"�iI8���D�>�����z��ֵŋ��xz�s�\���Ms��ΗB[4u�g�X��jY�ji��i���E$�$�qI4 $�q'є+�wN&Wn�c��"�o I�m�-��I4��� ՘�V�:�Ǻ�|DRM"I' RM"I'=0LŻ�n�����i�x���D�N���H@�$��K�o���!�܃SOkO^�")&��J���EV�"I'>@��R����if;`ږ~M�]��nܳ�i��uEt�l��ֶ�z��]�f1����&Wn�c��"�o�H�I�E$�?���Vb����m�I4��N")&�$���`��w*�+CZ���H���E$�� ���"�n���>�̃OkO^��D V�"�o�H�I�|�Fx+�7JL������E��#�)md[m�d���jk(]dF��pg���~~.��N,"�x�h&��ά�-�\������:�[���6\�۪̮��i+�L]�.�.���I�[0[YW]U�t��j�ݍY��ã4�$�q�۬e�g�e�Q��붣�ն���ˌF ����xM�i9�pVm!����]�F2�����Me��E���vn��lvm�5���l�ɔ+�N�v7Y����GF�!����
j4�vM�3<`�g�3��S���i7v�wZ�A�F٣�R ܏���-;=v�&�Y�,ݶŶ�`���9�#���e�X�So��edI$�d���P�x����3w|���56�9�"�o$��$��2< �����14��=z�$dI$�d��$���������&Wo>}�̋m��2$�q"I����1f��e�X�So��FD���d��$���}�v��x3���Z�-�b���G��f�8��g�hV�ѮQqͨ�u�yFn�Z���}���m���FD�N� E��?�M��F&�C5��_'�ݽ��2��`�h���'e��r�]h����n���;v�dI$�>}�3�\�Rev��ۼȶ���#"I'�H���F(34fk/Ǻ��")&�$���I�I$�,`�͸�i�����m�������m���FG�߰G���V����V���.Q@'������[�s]�
6]�.�Xй�i�`cI�����$��$��:H(m�G�x/`�ғ+��>��E�^!m��m��1A$����35��c�M��YI8�   dI$�=�3wjo4chh����{���mdI$�d����u-Pji43Zz��2HȒI��#"I'O{�����d���U�<pp$�ħ]�=��q���=�Ӥ$)c6�� n[I�����_�ϟn�#�����#"I'$�����b�3Ff��X�So��FD�NII8��1n��э��_oo2-��2HȒI��##�?~�Z���x3Zz��!m��m��0?�� �! ���S�����s��]�يuS���V:}�m'ܝ   �H/Y��X��\�Rev��ۼȶ���#"I'$����	�f��'�V7j�\ky���,]n[�����
b�u��Z]���JItM&�������D�NI�$�����z�qn�5�CF���d[m�d��$���F?�G�C�1t-������FG߿~��FIKx��~��Wn��]�����E��"L��I�I�a����1f��a4���&I�I$�$�0�$�Fҭ~X�NU3�.��6�V�\���ڶ6��H�D��aD擟`�tn�Ǭ�
��ض�Qd��5��V:M��ŷVIu�wi���eF�ܝ�v��Y9n�N��EƗs\�m�m��a���n���[4
�9�(��a:Yzu���]K͛c�z;t�Dm�nD��V���ڃ&7���^w2$��eQ���Θ��v�۝�8�lSC<C]-Kyymr`$Y��k�2�cRa����%]8�Fn��e�*��ix����n��7Sv��"����'ӗu�k���ֺ66SGcR:4so�j��6��x��a�x�2L"I'&I�p���KT�O6�|D�&$���2L"I' #��Yགྷ7Jx�������=�{�D�&B�on[�O�Ś�	&3wSo�� B�-�-��d�D�N#�}��r�ѣ[CF����x��{��-�$�qd�D�3�n�a��y��u�5�2��5�L�g\���J��t���X4ꜥ�ڽ׮=�Ʀ��=z��2L"I'&I�I$�>|�<���<Av�vwoa�x1���f�$vK���߹��O������$��I%�,�,зXI1���|E�n$���$�$�q��Ż�^��{ϰ�m�G��m�-��d�G~�Ϲ<	�z�|D�&$���$�$�q�@���ר<c��ēmC?&��û��'t�K���s�t�[r�y���Ԛ�S�n�gv�e���$�$�qd�G��Ś�	&3w^7�I�`�$m���D�N�����s��h�����}�z���$�0���Jw&-KL�4
�q��6��m��\:��ù�ԗB�'m��/��p��ϻ�x��=z��2L"I'&I�I$�>O�<�C7Jx����ݽ�[m�$�0�$�D�&���Q���a������RWMt��c��'<���d�.�)��y���{-�k�u6��2L"I'&I�I$�-f-ܺ�h�����}�[m��Q�-�-��d�G>���A�{�^���"L��d�D�&$����,�U�)����v�m���>�"I'A �$$���D�h�f���I��խ�d�G�[��-�$�qb�2o�u<	q=�w�m2�ݎ��XV�N,/ Pҭ+�E�6�C;�uf�z4khh�����x�2L"I'&I�p��ȱA�{�^���"I�$���lDI$�?�E�*�n��1fww���x�&�D�N"I���}��љ�$�ǻ��$؈�d�D�b"I'h�n��kF���o{�m���$�$�q}؈C�/�~���E��N1p���92����;�˷�n2����A�i4�)<;���s�O��7 4�55���q�5����3�MˋG3�x:p�����d�Bb�L�(�PB9G1�ܚf��w�̡�!t5�+$2�B�TȀ���W�sTNL��'�6kl��ֱ�w�t���[�S;��1^�jt��["��4>��3r>x~d�_��?9��A �y�~5pۙ��\jo�:}�S1���ݾ]�m]������>���5r����n1�CZ�ֹ��l�vkl��39�R\���������߇�.�1  :^����֕e���c��#E�,�۲5N�nR�lɖ\-����Rz22��=���*�%+uW:�V�gQ`gn�-��C�M���K��V��{W.��ݑ27L$ZM�i�I�h��ʽZݥq����<x�P4sM�-�		щѐ��H"t��v  f� $�uZ��
� c;Uucn�d���Ҏ�ݞ�����퓀��L�t�']qPj9�vN�h1��j�3ͶC)Й�4�k^�����&����d���Vfq��;\�uZ��X��;nŶ��ћ���u��@F� ���n�Uˠ�J��Kf�6��ۤ�oM��s� � s�K�8��f��m�$�u���Bc�t��7mRgV�z����
��O;c2��$!J"]����ڠ��v�Rܱ��P�3��Z|F^yўCs�8<X���=��e9%���� $������&Y�a5֎�z.{��0��<��W=�9�I�l[���z+lO=v3���9��v�GM��WQU�=,0q˥���� ۋX�J��^����zø-���mȅ�m�C����F��!*���ʽ@�v�<�l�1�mSg�1$^:��p�b;qs����0r>o6r� ��]�;y0峵��f�'Ig39fv����5�X��ƪ(�ʁG7N�Ǉ�k�LN�Ne�K���I�1����X1��m&��n���;�7wD]Z]Xl�u�5����ܳ�l�iјS�*��1LF9�UJKU�ObE���-v�R��X  ��;^ٶ��z��b���pl��Aa6�n�M�Б�t��V g���r�/M�S-��ہc��5�(8�I�Z�5����Y�a,��lN5�,��+�יj�t9���v��U�]�l�L�T�cR�U�s5+,�]��xr��ֹ�p�z]n5�wn�#V��%yIJU�ɀ`��n�$�NT��KV�6��m����m��m��_I����$�=��q�O�^B^HԮ�_)��{ʸ?�����]s�(S##�Zv��]:'�x�ɛ2�確9�@]�m�Lg'�erdt7>y8�*�94^p퍭��9H8�nc�w#��a5;��Dh��l���9�c� �6n]���\�Z�Kۦ�H��b���F�^����r�g�ó��+,[���ݚJ�:t6\C�1�*��n��մ^\�8��j���(A��;f�[�n�����I��0�=�g~�:�U�\+����
k\ �b��C;�v���s�n�˵�4.jFk.���k[�}��j"I'$؈�I�|�T���ř��>D[m�$�I8�&�< (ϖ74fk	&1�����n�D�N"I�>�8�Q"�ݺ�h��ѭ�w"-��~͈�$��lD��gՊx��=���&�B2I?��lDO�N#� H������4�<fE0e�Cr��d�����������1�v֎�s5cI�����Y����"=�{�D�b"I'xB۵>Xh�љ�'������߿_�L�d�0��J���^>H�Er��:w��؈�I�{�ݸ�ѭ��^'܈���I6"$�qM��|X�1�X�n�ַ�I6"$�qM�	 +m�D�g��������>D[m�$�I8�&�GϨ(>�ֆ`h6j�7�Y�#cO77(ͲY��77Y�6�Zh���������n��k�w������I�I6"$�q�ݹ�h��ѯ�D[m�$�I8�&�G>,
d�,z7Zk[�$�I8�� �H�(� ���D[��#�ߣ<�C7CY�wwvc��/{��mڈ�I�R��DO��4nk	�f=[��$؈�I�I#I'����#pGM���Q.��U����R\�#Y���g��d6�������5��
�m�D�0d�qH��őfd%�F����$g��(�m�-��$������%P���`���ݙ���"I �-������>����u�����o��m�m�D�20�� 
�H,�I� } ӶN#�J�n��4chho1��o�@6���m�'��������̿�kK5]]�̕����\�ɰ��z������S��S����1��Z�ka�o��F�N"I2I8��~��U�f��ٝ��m���k�o$���雛�wXy�1�����$`�$�$��$����"�u��CCy��/{��m�$� ����)�sq
K^�l5��H��I�I#I'�` ]�@$$�Sr��i�����4�D��
��" �b"��s9S��&�CF��|`@��_��ef��%m�suwS��@�R�s3���uv�B6 �خ��ӯjys�m��Ǻ�uZ���;d�r��cG��c2S*E��6�Ӣ[�v�������J�p�޻WJ������H�=I��^��<��9�z�U�e@cl�t��
�����œ��A�CKNZi�5����3�62���;:6���n6���g��;5Mi�z�'�ۻ�ZHѱ]�v�7�v<��s���Y�[���֣l�^{��`�v�
�3���;����$�$�������a�����<Ř�n�|D�0d�qH��IAj���4chho1�����I#I'$����@�Z�ki5��H��I�I##Ā���A�K�f�k0`������o$�$�D��0~�t,�����6�lɮ�);e�z9�ͬ�tzu��s�T�r�y�z�����a�,ǫs[�$��$���F�N"��f��Z1�47����?;��f����湕���Ӈծ��l�n�t]]Uƪ�:�8����[�E�ON�﫪��:���4�d A$(�0  0�����K8�$gĀ���MYCAk���{�����IƐA �m�m�G��3�T3t5��v�p��m���lDI$�$�?��7wswXy�1�����&�D�N"I�$���蛹w[��з7F7�4��)pv[fЕF�,�
�J���r���G<��S�
n�cCF���"�o$؈�I�I#�/��@�Z�u���$��$���F�N#�}R�f�k3����xm�D�00}JD0�!�u�ήC����c�p�[mP4��H�:N�'�+������a�,ǫs[�?�
�X6�x�$`�$�>����n�c3Xa��xm�D�0d�qH�����E���z�V��,�Z77Oe�c���H֘юڹ#¶��α����v�2i%�7XOq�"I2I8�$c���o���K�f�k3����xm�> �Di��6��������~�����<Ř�Ǎ�#��2I8�  !m�m�G�QU���f6�m���o$�$�� �0�A�F�9�>�>��6�Z�q�����#"I'$��$�G߿D��懩��	��wVbѶ��
�n����\u]�����$v�3n��j�f�k3��滛"�o$��$��2?���7wswXy�1�Ǻ�$��$��2$�qm]����c0�s�ȶ���#"I'$�����k�i-���I�o��FD�NII8���eJ�����K����l�m��2$�����ۅ ���n�k�6��� �[x�<ک]�F�#��t=[ͫm�g��+�E�7�i����pq�6q�G2J#�mV�"1vieݴ�j�G\]u��sm���T��.:�v��tj�콊��`���������6��f����1�'n��WG	��7cl�DS����k�>�ca�uC"�9��X�j#q�%3��b�Cu\�iDwnK�un��6Y[��˺�������y5�;ef�J�oj�\F�.nQ-rt�n�qI7%^�]-��z%y"OsC����a�,ǯ���g�ȒI��#"I'�*�v浣q��o���-��2HȒI�}RM�F�}�q�Ao^4��|EV�"I'�H�I�}�<�C7CY��owk�zE��")&�$���I�|��D����$�=x���E$�$�qI4�$�G��Eթ�����Þ����Q.��U�Zzv��e�.�����v��M#���kF��kF�1�y�i�x���D�N")&�?�>��Z6�Ɠz��F � �  A8� 4����*�iI8xQ�b伆`i�%����^��{��"�iI8���G���Mћ���I�׏[|DRM"I'�H�I�_��7nkZ7i�{ϻH���x���"�o�H�9K�EL�][ú�K�vm�̯eΆ�JD]S���g��;r̽n�ҵ-z��[t�$�DRM"I'���fT3O1.�����m�DRM"I'�G�(��`��775��ǯ�|EV�"O�q��@f��D��"~u�&i��t�6>뽚�f�m^z;���񩦳l����/?p{1�T�g
{�78���l��ՙ{��j��j�����������M*�嵵�6i�kKr�[��<��|�_l�-��7����s��q���l5���ڮF����o��-�ڱ�m�x�޸G#NL�
����h�¸.
*D�\̘�"a�^%�p���;��xnf�q�,9+00#�g:6I�)*-){�a��ι��_ywS��_$q+�|�x�*��V��^���"�}Q5$>�}#�z�{S��>NS�J54C_��~�8��U��kF�0���[m�"�iI8���D�}����{�����H�I�E$�$���w���m�����;=�d�P�|��h��2�B�M%���6�R[���-���Y4�u$5��]�ݯ���x���D�N")&���>��7swXM`x���E$�'�'�H�I�_�Q�n�ִ&7Co�="�o�H�I�E$�'�A|���z�5-ׯ��I�I$�"�h!
R|XNd�,ds��į�O���|�T����1v�v�פ[-�<$ܶ��x���)%�	u,zn��QF��&���׳��ts�5�>"v�h܁�'<��j�^Q[������ۤI$�$��$���Ш�7nkZ���xm�<F�X6�x�$`ϡ����A��Էq�"I2I8�$`�$�?�A�J��x�k�����m�$��'�8�$`�� ��w7u���=|D�0d�qH��I�#�|	B~O�ſ�2]��%�[�l�q�ہ�s��t閉k��ızN�H-�i*D��qK���p�]5�Y5;d��v2KR�����Xϱ��dO-��1���\r�l3��Uu!��*��~6O�kt��y8bh������Ƿ5���� �FMո
lMB}ra�k�i��A�`d�F6z�(�z�EYp��6`��!t�+x7gG7�q�٪y��?a����u;F�c��-�궻&��Fd�.9��J�0�* �k<��'c�����`3ޗ��F�N"I3�C����Hf��Kwu�H��I�I#I'���T3Ob�}���m�D�0d�qH���A7F�n�	�'�=|D�0d�qH��I�_���zƌ��{��m�$��$����߿i��ߏ�we���������ײ��`�v,e�R�TF�vݛK+u�ܳMIB�DwkC�зs_$�$�D�1��o��伆`i��]��{m�����`��6k!�Ѱg��qHψG��E����&�<x���-��$���Jl`�$�=�P��V�h�a��׼G�!{����m`�$�4�$�� �}Պ�{��k�$��$���F�N"|}^-��:�nڡ^]-������g�QX�c��7���3��M��Ř�_v�>�o$�$��(m`��h�swXO0'�=|D�3I ���"�X2I8P ��<.n�ѣ1��o^�>����'�߿vus�,�)��@đ�q��
��s	%��p-���x�����"I�@V�x��h�%�3if.�ݽ�����I#I'$� ?���Yq���Kǫw"��k�����N�g��#r1v�X�5c1׭����y��'�Ǐ��-��$���F(  -���������zz������ J6�����I#�B����If��Kwu�H��I�I#I'��	�K���v���|��"I2I�ÿf��--�cS�T�'0~�O�0d��a<��<x��H��I�I#I'�%V�x�M������ʺ�z��X�튋�h�u�t,[M��M
k�cpn�oF���o[�m��H��I�I#�B����K3^n%����$`�$�$��$����ږ!��}���m�D�0d�qH���A��3u��fkO�"I2I8�$dxB���}�`��Ѹ0�kz�m���F�N"I>?�$
#�v�cq��r�/g���f�R�+հ�m���G�v��C�����1�a�K75�[����c���	5c� ��0�J�Ě�zۭ�s�Z\l;�*�鍋�΄�c���E���n(n�vńv�m��s�y���]�c��v���0��+#�[Y�;u���Mݖ��F�6�1�֖+s��N�F=g�[h�U�,x15���ë�t=������)@-�v�ܳgcAu���=�3�8�^+<�3��;g��ǈ��#���G��0|@�����N#��%�f�Ļ_v�>�o$�$�D�0~|�V��[�<����ǯ��F�N"I2I8��}�wkz7z��o[�m��H��I�I#�C��f�%��n�����$`�$�$��$���f%����wYV��H��6t�$���0ݎz;7O]� M��;�m���Y4۫Ctb��9y�����I�0d�w�@[k��un�ź����<z��$fB$�R �� B�H�~�@�ֻ�_�kI'������'����_m���F�B�om���zIcou-���I#I'$�$�GϐM�X�`l,K��o=�m��H��I�I�b#����v���֩�d�"����l���v��T�4nx��[�ϵY��g�_$؈�I�I6(<' ��G�&n�k�Ԟ�����"I~g߸G����$�?�dm�a$��Էw_&I�I$�_�.Ԉ%(��%����l��L���x�9���G��&Ա��v�ů��m�D�&$��� ���p��mշb׏,�i���I�aI8�2L"I'�߿�[�3`�lwf���f�*t��̓��x݅QhV���Y��{nV�������m�D�&$���$�?�?dz�0�m�Էw_&I�I$�$�0��I�}�V�`��1��o<Z����I6#�P���[v�>��5D�n��1f6��|D�b"I'$؀Ѵ ���̣/܇9���ю\)���e8˘��F��S���.�m��qG��?�<��.nկ3Rz��m��E��"I�$���lD|�� �������[�35jWq]�3�//f�jd[�N&�џ*��y.��>�u�zI�o[����lDI$�$��-�G�E�K0`Ƙ�K��&�m���lDI$�$�?�3pn��f,����$؈�I�I6"$�q`���m�k4,m��|�[x�&�D�N���Q��[z5�Y���խ�M��$�D�b"I'�w�AH$�i�j�|�͛6����L�;���d�-Nli��LB���r�����6#�E�Z�;�v���Mn���ǜ�Vs����ئ.����H4�E˝k�<k�5ŷ��#�om�#ٺ�cz[Uގ���!#1�#��}���A`p���]N�뭯<wu������|��fG9j]⻎��'�m���+�u_Y�歬�5���\��	L��Z���Ϸvn�������Y�L�"�;]-���'��E�
8�K S��ڍn�l�����ca�?hP����RaV��
'N���M�;!�py�B�vzu����Bm���Ys�Kbql�`K�ʝ^эV7\��pYFy�Q�J�Q�US�[m��Hݶ��� ��@ �>����id�9ov�9z
�;�ݶ�s˛K׈�n���nݻb�����!ݩ�u�i-�!�63���^�W9ڥ��86���,۲��Z�a�	�U{g��F��T��E3�&�B��t��s�/P�е( [@-�sm�ww[I�l���$7F��4��ƨG��w���m
kU�;Z�[��l����I��7M#*�\8n��s9�}���ī�ɹ�-�M�l�wf�2�JN��6��
6�M[%h��n�#��l���3�q�UM���ڳ��pV.�$�[�͌Y�j�6��Vހ�8�8�0�q�Z՜��sn��Zy����+*Nƺ�F��b��|�v�mOvv���k�s6�w�e�s��N4�;H���T�D&�.��Ŧ���km�T�7g�:�m�X�]�ʄ����ڵ��#Zo�}������F���#+b�%)b��&w6�2��UC�>y6kl��Ǘ:,��I�`r�u�6�z�����j23UU�*�.w\܏vQ�����c1�mK���<>3Ŏ�h�=X�;�VZ�Ul	lM�mS�%'f���m����NCK�N��s�)��S��hy 5������l�J�=-�j�B���lv�W ���m��읺���m�������8��U竸)z��J�P۶qa�8�%i�y9U����ɶ��6�`Ҵv�;-ƥ
r.؆�w�	��"g�m�
�]���^��\*}�W��툎��#�64�+6�R"e�f�eP!�-�Kԋ`t�<�
�f���tquR��K�#AYF���,�#ss����Ѷ�U�)/��z�
��n�����7�WJV�6.E�+�W�='j;���D�����?\3�C004�0;��d���³d�ݱpouR��ce.���2C���T�g��)c^�p\�{s�',�DՅm���x[c��cl�Y�%lv-$[��r�ۡ��D��!��Z\��k��A�۲��HO^՚�ͤ]�[K�2䆶h�+*i�1�Q 1f�8޺g�q��ɷkgJtF*����a��ϧ2<�+Z^ȃ�8)��]�������hog'3��.��.g���ô�{�i����݁{/$h�G������9L�F���n������Y�4�b_��&�}�x�&�D�N"I���A�7��b�m7��M��$�D�b"I'�����ƳB��m��m���lDI$�$����Xŏ[L&��"L��I�I�aI8��Z�f��v�ů��m�D�&$���$�;��Jn�^)��<�oj�\kt��nU;f���vq�#�T���#��n�<Br�@`�M}���?&$���$��@ ��"P�g�}��hX�����m�FL��I�I�`��Sm��c���Bk[�-�p�$�D�&'�8��z�H!�1��o<Z� ���{��-�$�p[���.n��Ř�m��I�aI8�2L"I'���U�c�ƶ�Yś�3���c�0�����-���k-,����.��7FH�^cY�cl6�s�-��d�D�N"L��g٭��1=�֤��I�aI8��$�$�p� �~J��06%��f��=�{�D�&�H@$ID\+�w��df�5u�WXe���M�M���8�����j�s��l�ѱ��f��]J�󻜸陌��:���v �'�u�{��>�#����7�a����ֶ�&I�I$�>�&�$�������ƳB��m�s�-���r[�[m�"�i����7�����f��a U�幣s��ݗam�!t=P�fӌ�s��x<3K[�z�K3[�"�iI8���Im�G��� ��Ļy��"�oF�n�m���I�}��rf��7�������"�iI8���D�N#�+����k5,oCo�="�o�H�����ڷ��L`��S���?�H�d�޵�1,lbY���H��o�[t�$�E�����a�v]�=�H�#D�v}���lsѵWN& M�s����=�,��i ���v��{�G��{��I�I$�"�i�ܙ�7C�ff6������D�N")&�$���
���ףt,oCo�="�o�O�!m���-�:�n�k0bX�ĳ5�"I�$���lDI$�?���0�X�7�n>D[m�$�I8�&�G���h͘+���{Nzŵ��m�%K�.ç[��*�V�WFh�˸[vI��+�c��3��:�ny���&��Y����H��b��6�t��;t�sd�׷<cKg6�W�^k��-iK!�K�6h��-XU&��[#s� �ݍLtq�Z`��)׸aS[��ž�a�t�y�)5r�3F�i�L'E�(	s%��-i�������V������6�kQGd���	�'��㣞xd�9)xų�ak�u�y���������������$�qd������}����ƳR��6����x�2L"I'$؈�gٺ����cc����&�D�N"I�$����ei ����y���E��"I�$����mڈ���WP�kř���m�M��@6���-�$��s}��/���W.ђ����7u�F��sXFh�r���l�⋖�p	�Ϻ���V�n{֛{�e���lDI$�'ܓ�g٭�[��y�fk|D�&	4��B ��H C6��E_,�$�q�dU�����ۼ���"�o�O�I-�*�����SP�kř��{��I4�$�D_d�>�' C�{v���Z{�ޑm���$�n�m���I�t�>����mn�չ�1�Wp�d�Qym�֤ӫ�$W7Vϕl/^���ϭ����kpbY�0-���H�I�E$�$�q� �� �k���^>�-��I4�$�DRM#��ϸ���׋31��[�'ܓ�I��H I�đ�8 I����8��!�.�x�3^��;�m���$�$�qd�G�f��nb[�`M�7�I�a$[m�"ܷ�I�R }�e�t<x�i6�^óoA'��ݟ\Xɖ�W��`@�{�+m�!�7������a����2L"I'&I�O�qMZ�1�fci��I�aI8�2L#�q"}���h�z���xD��"L��I�I�a���'������x��I%[��������?~��U���3S6�@�H��w:��P��q40��m��"�o&I�I$�$�0�>X�'��Ø�)q��Tn�e�ur��q���tV���������zݤT��.�V�o��r�"I'&I�RJ���}�!=���!�5�Os���x�2L"I'&I�wς(��Y��X73|D�&$���$�$�q�`V��!�����{�E��"L��d�D�&?�}�5�ΰ�1��[�$�0� H���E�n$���4� �Fhz޽[�s$н�Kr�Y���v:�p\�]��u4�l����5K�f�];����7ۛ�d�(��[�g[K�˴�͡�G��#��l��d�m�V���u��c�\��2��b�K5+�]]��8]�e nXC{b�IIF�t������k�8�m�/9���:�Rəv6�z��4��ͫ��t�5dܲ)K��}[.e�q0>㎆�[,f�T���}�C3%7��mt�vKxUS����)�9d;;c4F�X��������d[K71�0=[�Z{�y���x�2L"I'&I�wς(��Y�֐�ǭ�d�D�N"L��I��!R���p ��{��{�G��{��$�$�qd�D���&n�ΰ�1��[�$�0�$�DRM"I'��J\ś�ո���y�>�o$��$��20|�m��1��Ys$�S��s��Zݟi�u��kg��N�­�i]f�d��T��w�~�����߿x�~�>������+r������2-��HC�@
@���hC�#	 �[~2,�g$�xQ�%˛�t3�,�m<m�6�ȒI��#"I'�E3۫7F�q�O��`xB���p6�ȒI��##��E�Z������f���#"�����D�~��*���E��M�g61r����ц5:�%�6��۪P��Yf��a.�z��"�o$��$��#"}�3pn�u������Id���FD�N#��&ׯ7Z��S֟c�ȶ���#(O�PJ�\x�!/��5��'QS���^a��(�?3��z�w+��"E�#�̻x"8&&Iu^�.H�e�7٬��΍��O��\i�E��\�@G�3��J�dL��b��tE�p��D�E�<�	0p��*��y:xn����kɭkV6W���q�6w.9���r\=�82��]�V�{s^7��농��ij�Lj���l�Z�yN�{�3C��k��s0%�9�4��j(�0v�q��&f!,�|.���+�yf�s�t�9ώj��=�i���ju�k�w=<���R���������т~�ᩁG�l�aB�ˏ�f`(YD~���E!$1:�f=\\/�e���������-cr���{��i��]{��O�T��Sگ�9�#s�s
ގT�蹊7Y�䛫��,��U���ן=��-dt�"��Z�ķXI��o��FG�$�d��$����ʷha.�{�y�m���$dI$�d��?�ɡfŭ:��vk�b0�&�M��ҋk�!�Is;i����p�I�8]}�!9z�v�U�{����"I'�H��x���5�u<ֳ��d[m�d��>����FG}Lǭfb[�$�5���#"I'$��>��H�u�%��u�2-��2H�����O�Q`���(�% `��q��Z_��:��?ϵ@� $O�ȟ=외7C:����z�$��$��2$�q ������u����Ӷ�E���c�i�a�qhEqE��@��y�]�KL4t�?����{��d��$��@�E��?��U�z�f%��O1��$dI$�d��$����/�q�%۸��E��II8$dO�rf���3O[|�2$�p2HȒI�|��ͯ^kx�y��-|ȶ���#"I'$��p��?�YZi���d���g��l�m�Ӆ�v�F:r�om. ���Ʀ��p^�x��v��rݖ����7(A�l�v�ڡ;v��`r�st�FN]�T��=Y7���n�TS��	N�1)['7u��+q�b����÷�+�ɭ�c�h��p�l)�lV�mt�ĝ��:�܅�;rU�S��W(x�-�Ke���ݫivjLfN�C�N!�+w�6U�����w���w��5��l)�g��c$���0�jHJ�b'���9�ע����{]h&�lMby������I8$dI$�>}K��A��]��[d[m�d��$���F?�%�L��7C:������m��$��2$�q>/�|�淘��z��̋m��2$�p2H���>L�7Z�ĳZ��o��FD�NII��wߏ��I�f��[�lRV��a'O#��nό�O2�*��ɫ$��$u���4�SB]��[d[m�d��'�;��D[k"��2����6���$a �<�CJŬV�K����="> <�6�����k"I'���7�ך�b{��{�_2-���O��x�n�Gϟ&	����%�<ǘ��"I�$���lDI$�'Ծ�e�C40�7q�h�m�D�b"I'$؈��A�.�^^c<%�Zlu;r���T�ב㫳B�g��n��q�����-\���M}���b"I'$؈�I�O����涱���{�{��x�&�D�N#�ܓ����3q��K41����I�$�8�_�i��Ɯ��/�k�U���ڈ�g��|��ˈ ��avn���%��M��$����D|��nT�Ӭ,X�ou�M��$�G�6"$�q�������su0�쪧�D��"�r=r��ϳ7J�z�{�<�v��z�+c�]=h{܈���|�b"I'$؈���`���f%���y�u�M�x����"۵$����}�ˈ ��avn���-��M��$�D�b#��/��CcN��1����$�I8�&�>A��i�NtގU?��C$�~�����,S.��m�7S���D[m�$�I8�&�G}� oqkd4*W,�]�ã7+]�����#s��wC�l�[8b9�t%��u�����ɱ$���lDI$�?�_hˈ ��c;7S���x�&�D�N"I����١��ZY�^7���&�D�N?�([v�-��������`cu=q>��{����n�D�N"I�����3q��u1���u�M��$�D�b"I?s�{��_���7c�d�-�� �5�L�ıKT���`	�vٶɸن�-�L������%�jGA�x�vz�v�U{E�c��Ю�m;K�L��N-vK!��Ŝ����u3��[��j�h�}�����Sj�ۣ��)����n�X;=�9-�.F̑GD�c��N�XZ݀{������!�.h7Hgt���":����N�����Z����V�_�����L��U�:l�ٶ�D�9ۿ����������0���h"� g�cW[�{��j�tc�CF�����h��~��I6"$�qH����l��ӭ,ǯ�|D�0d�qH��I�|_r��m�4�Sя1��o$�$�D�0~|�&n<�An�Y���_�%[k�o>H��I�|��� ��c;7q�l��H��I�I#}&������x��F��f���$�hݔ�Zb[�n�n�wd��Xǟ[���4�K�י���F�N"I2I8��L��y�-��c�o�������xO� ���o߶�H���}�3q�b[�����|D�0d�qH��I�}�����n�f���G�����[+I'$��R��cN4��y���$`�A6�����N#�����V�/<�Kv]�X�.�^KF�St�-�aB����4� }�v��UOc[�����I#I'�$`��>̙��1�X�Vfk�$��$���F�$�>����$�.���X2�x�$a��L�ƙ�kFb��~ ���_���_���}K��i�8��z��k�$��$���FG⬖�%f{i�f�z1���"�o�H�I�E$�>�|v<ֳ�5�֖f�6�ۗJ<���'Z��2Ǌ1s�F[nֺ����\E��f`M��5b�|DRM"I'�H�I�_�R�2�	������-���F/�4�$�DRM$#�D��i�8��z���Um�$�qI4�$�D�}^˭��3u=��s������I4�$�S��0$Y٣QD"�l-D���3n�6������ $0�	�$����#�}�7�ěk5�u�I4�$�DRM"I'����Į��^��-m���f�m�'��>�>ʥq�5)Ǜ`O'X�!�havn��zE��")&�$���I�|��/�07�ZY�^5�����?���Um�$�p�@ڔ^�n��Fn����}�{������D�N")&���}�3q�n�M��֭��x�U�H���E$�)$�����f{3؂C40�7F�"�o Hn�n�m����Ϟ���zq�k�P?J�߹"�I��Y�B�bqʈ�y�J��)�"�o�ES�/�~Y��"ب�U�~�Y�������~W��_o���_�����w�������}���_���U�o����?��ʠ������_���� r� ��j�]��_U�ww_Z�����ݟ�7_w��~�k6/o��|�
���%�"XT�%�L"5,��hf�43Q�22�524VFB��RhjQ����hj22dj�2hbdh��F��+#J�E��hh42�2�2�0�ѡ���Q��VF�25Y���M�245Z�F#��MS#KY`ƣ1-���Yhl�hcCZ�F�`Й�J�ʲ4�cQ�hkCV���Z�dd`���`Ԛ������5#CJ�š�����2��Ԗ*�@��LF����V�Q��d5,�VCCG�8L24�C##�PҚ�#RZ�D�1CP�CK#,�,�5Z��!�#MCSCL�&F�P�25FCJhj��2SCE�d����k#b1���1hd�40`�b��#PԚ�CPԴ0�CTd4�F�d5R�hS!��J���²FC�4X2�C&��j��K����j2�F!���j��2U��5&C��j&���b��,��C&����d11����jSP�L�Dj��`V%�d0j�K#!���j-LF,��%��2bZ�M%�d11dZb2ĵ����%�CM%�!��dĲL���XX���d�KI`Ĵ����j-F%�İ�dȰĴi,1-LKSҲ�E��,K(�,K�JUU�e����~*���:8��9{�p�O"�^���m���w\??}�ol�.�b��X���׏�� 6�T ��z�^|wĠ��ڐ��f����p���ٿVx]YᎼ1mp�J c������z� <�1��~~}8q��,���ofP���� y�;^V�Ž�q��og��~�}|�y�9��7>�� 7�c�]�����m��ۮ���@e��
������|~�����z_��1AY&SYƧ�X�߀rYg��?�������`q����������R�J �*������		 ))'�p|P�< �;�@^�:���<�&��� ��  /cE�s� nx��nn�h(��=��QD��ܡAﳡE�ۧ���n�|�\=6�� ��z^ګ�;��+�\t���3��
��w)T�7<@Un�s�J]��R�{�]^>޼�s�+���_7<@��ꮰ��ܵ�w7K^4�㎩kwWum�>>� �  � 4ړ#EJPё����`�d`�)��T�h�T �  2h�   E?b�HҠh4       �E��� �  �0@  � �A�ё=4��M'�i��Q���B� �Jh&&�&0 �0#�1�v��$	��s@T@�(u�y E6�@M�
���  �Q�?����n (�cY0������~��~����&��{�o�������|h��&=�}�m���7BD���PQ'
�h�Cz�� ���N( (̊WY���I&�]��Q:iBr$6�-��XF� Q�X�Z�%���W��O<��o}��)��}U������*�
 n ܈�Pp��@� 7" n�p��� �@7
����@@Ց�qn���o����*r'qP���T�t�G���9�[��}���{]�M����&�h�f���7Zb�1k)�F�b�E����n3~Gf��j@����h��fã�8�9^:w����x�K2]y�Vޥ	�7�\O#L��\d��n4]��ť�Ȗ�t��U�-�4��	�V�sp�dk�6F�:z8���ʨ
#��:���hF���\��vo;-��LX[��&��tR�Ѫ&��vi�p�hcS�ƠG�.h�Q�+�kڱ'��4��ڭ;��v�%�6�Ť�t����Ʉ��u%,I��4F�X���oy�XǈJ���ԛ��k�����gG�uRd��DNpX�ɚ�H��*���
�bu��af�4dU����j��8�`N�kD�&��F��zE�?tii���½�qkAx������٪��L����2gdmh���t��!���,���d{��I
5]HHN���7�bk�7wѥ��`��l��f�Τ$��H���<�:����n�"[�V�@�����۰U1�&*'�[Z�3#S�)$Ãz5��	�5�`����5�ɯ'��/!Q}�KZiֲ��wz\�uцr�Y�FBN1!��5�u���Ձ�Z�bi�C)��9E��$��11��E�p3Z7j6Do}q�'}Fp,�B9��Vc�-��i�E�Sh,��!7f	�LnW�@b��d��8��~u�]o�z��(��i$Ƥ��ye҉T�,H^��k-�R���mS�D�#�߫�m�y�8a۾�x����l�"�2�o��n4os�kx�_v�O	Kq���o��y�eN?Cʼ�ܕ��.k�m-�Ȫ{�^4ӕkmK���������ҭ	a���s��6��h�խ)�x�w˳B�41Zރ"�3R�!�).m�Ǚ���+St@gl5�����X��K�8u���=���,5$�u�ܑ+��!i�q֩SlH��Դ����z��6W�u�EX��cq�K�sx�h����3;��+�JJ��;��jl�fu�9�y�Ί�Дy2Ti����Z�f�39����`h�\b#\�p�h��3l�LM�5�^��O=����U����8�rl��ǧ���g�@@F<��sr�ˋ� �b�!!�@`A���qtGg9�S�-����3Z�5�`�(��ÿ��$����.�y93[����gHX��89q:���n�W�ݣ�N�mVս�f��q�p7:��ͪE��N��k�����v�k������rmӘ��1�pe�Ԧ~}������i���}��ff�p����~{�h��Sg?�.�CSS �=�]�{w���������X,�Ui�����j�����av�d���V�3�bN8&� m��m�� �mmXn  #u�
F���WV]
U� 
|T
�
ګ�<��R���.qbj��`*�R8�t��׀\�m�&�;
).ҕf.���J؛�2U*��[$�p��������i�:��c�jc6n���9P�Z䩨m� 6�	�Ŵ��wYYzM�                           h          m��               �z        ���k�Nշ��l�3��n�ɫ���y���;�4�i��U��̪���UU8�Ej�ekv�*�X)ez��2���[*��U��j��4�۷nlB�n;2�J`	C�n�l�R*&7�Z�֔%������T�V��
U�^X�k������y��Aճ��Ax��j_��pō�vP*^Z��Z'Z-�6� �:t40u�gj�v��cvr�Gm����΍��֓m�r���ӷN]�Yۡͬ����5�ChV��i�<�ˋn5c/ӷ&�8Z�Cp)\�|�e����X��;t�.�7=��G� �um��77o4����м:����5����j���K�A�ljrfr�FEU�*��"�z�+���j��C .۶Z5��Vۑ�)UPAS��º�8U U�+J�l@�UUR��RR�X:�m�ɴ�]���zT�-��k�	ţ�A⑱ODd[N�T8f�UJ� �ʽ��
���VG!KvQ��� \�m��� ۿ'w��/�\�k�CV���6��~}{��ޅ��`�9��z�`��e�h�^\[ؗfl�6ط�  W�D�I�R�ol��^g���]��7\*��!P3�+V�g-�;�uV��՟ ��&m��M�n�}���
1UT<�qjkcH��R�[[N4��+V� ���]l���G�@B@��Ͷ�� *�U��
�Z�RZB��*�RUej66(ԫ�� ��Ͷ��kh�pa��H F��UR��r��1( q!+F���[�6ճQ��   �9�r@u��Rѭ�m5t�i���6Ƹ�r��u *� �ڷ��t�i$6��� -T��u\q�\eQ�8�B����i�]6Ih-���	 �l$  �����p  h 	  Xa�M�` p���O$��N�{;��t�N��k�Q�6m�h>���d5��#������ ���G~���b67��A����[�Á�iQ�AÜ���������/4	�
��S`/$Tp��K��	E%j� @���� ĸ0�x0""H (�^�8T:P�U!�<�� lW�	P�6��<�%>"����K(�4Y�1AQ� A'�	�NO@x�bv��+�'H'@���0yP�(t<gn��`�:|LxN�΍��~
$^<DA�N� �M�ZC�h��M�
l�SHb=��WgK��!'���<r �"��$j=���.�B�NS
��D��.)�0 =|�D@� �*����E����˴>A ��(J F��7��|��kx��+��Q���@�В���dy׎X�Z넛V�K��	�7׍^T�km�n�        �m  ��O,n۝Z�冭�t�%�"x��Я	�iڇ��nv�7)e�(\�e6k�!s��lv�(�+7;[�a˱k����FVx�[��	�I`6q�C�����knsJQ�+����7w# =����ۭl��[f�n��ʘ�ƹ�N��c�jzz�5+2�g]��>cV�1���R�Rۘ���e�����4]{K��[��U��ZX�8�K��
XT�	C!��7��0Z\ ��r7/�94|���۞z��#����
^rj����ȵ���[�[a�p�ѓvkQtx����K�&j}Ԗ�i,�k�;��!2��)�yH�s���|��~��n�w��,�5s���S�w2�+�r�5ț��[�,AHȍkQ�<�	���e[��\(m5������9(^w�kl����zRs��ۄ�P
��GJ)��f�竚����ؖa�&�ye)������-�{'e��7��������d�j&H��h	$���S{�H{�j7�쓼�c��o��w{@ ���9�XQ��ՕM�	8���o@=�&�8��
���n��n�Zq�֋6�-N\�pӘm]����%������ח\�cͲ��{�����܅Ы���ˉ/R̺�f�RF��-ѧe�U��lo�$ﮇ���)$�sZh k%s1M���R�L̅�ŎG7]�����Kd��y��k��Q���N#@�% ��S�$�rM�߾��+�2|�I�4]�ƊK�u&C������p<ɐ�!�t$�C"rYm%�B6�F<Zk2L�$�G~xk��L�$��V}/=�E'0��B��C�=�~��d�rL�˳�-d�C�d9']��^ev��Ub%��U-SK6�`���j
�����G�jMC�{����p<ɐ�'�g�Z�=�u&A֑4��2Oty�&�a�rL���u�W(�HVX�D�7�M`�d91w�2�\2d9&I����N!�2��0��p�I�rړ���nN!�28�Rw��Z�:��5r����	������jZ�42�զb����"�mь[vh�N�V���7Ǉy����������-�Xߏ��/_t��i��Q��ɸr:�vq隸���u&��V{�e�=��RdƤ�7�^�,��5��5�\��TT��,��28�d����V<Q��\�T����P�'���pܜC�d9'�o̼�̙I�yvyŬ��5jGw��[���-�ز�\(���y�!�2Oaߙ�+��I�r=}��r�\Rd�W��(S��{z��`6��?j�A�63$���Z�i�1�,��x3.�Ɠq(�Ɋ���'��٥���a¸���$�:�F|N�c,2с��&��k��h'�:Qخ���'�N('���v�I	�)����ryzuͬ�c��w&�ݩ3��{���G�2X<CQ�_Mu�E �vZ�[uɽ�Nd�58P�&��(J��`�%)BP��ǹ{�y��(J��(J��5�%	BP�%��(J��`�%	JP�燼�ˁ(J��9���(JՂP�-	Bk0J��(KV	BP�%)�o=��<�BP�	u`�%	BP����(JX`�%	@J��	�	�d&��(J�������J��(Ns�(J�W�bX5�`�%����n���IH٭l��{���]r%)BP�'Y�P�%	Bk0J��(Mf%	BP����(J�����P�%)Bs�%"Д%	��(J��5�%	BP�&��)P(J�׷��k�D�(J�����(JY�P�(%	��(J��5�%	BP�'��z�z�J�� �9���(JY�P�%	Bk0J��ZF`�%	BP��ǹ{�y��(J��(J���+�`�%	BP����(JY�P�%	By��uo�0�[�5���ۉˁĀu�wI6��*�r���Q/2,���;nH�quʬ�bt�t���v����瘪Kˉf��""K-���E�a���6r%	BP�'y�P�%	Jk��(JY�Д	KN��(J��5��?�(J��:��hJ��b�%	BP���(J��`��	BP�������J��(Ns�(J��%)I�!(M�	BP�%	�0J��(O|�ܽ�<�BP��	�%	BP�&��(JR��%	BP�����(J��<�y�	BP�%	�`�%	BP��H�тP�%	Jo0JR��(Ma�P��&�&�.����]�ZDB��,vG
�|pk�D�(J����(JY�P�%	Bk_�eL��(Jy�P�%	B{ƿ���(J��9�R��?w� �@r
Д%	�%	BR4&��(��%!�$	��%	��=e��J��(N��(J��5�%	H��!(L��(J��'���֓��Τ�9�P��߾5�uг�ȕ��X<\}ho�4�1�X�[&�*f�L��ji�-G�^��\N��9ulg�sӭ��������:�vjMÚ�;���3�w&I�]��=�=>և�9u����-(O��U-��)#�jkC��C�dt����y��#���~15<'?������rz�:��g�����ɨr�pb�Љ��ïz�/�¶�y�Q�/�O�z�ؙm%�7���@?��g\o�m懩2�Q:Q��?q���p��a�B,��Mˑ�� 0!#(���g�٨z� � �v�� @!���9���8����*;� s�w&I�69�?~��[�t�ԙ ^����;9rR���@�kf̍Ͱi��F)���^�6�3�:�7F7�V��Cu�Z���%��đ�u7j�l���W-�3N�m��Y!��J<]w�d��iO�ZiMG�^��n��m`�w�t�i��iPQ����Q��x��x���+�e�R�-a���{8֤��!�=�~��cb��w&��|��g<�֤��cP�����p1Ԛ�#�ۙ'�kQ��'M�5A�+����F�b$�`��W5�h{��g!���ԟ�g�m�Q����08�p�h�~��~3��L�G������MA�{o�z��0�L�$������y�ϼ?;�ͼC�/���J�,��Up�Y5����I�9&C�g���8c��8�ɑ��-�}�I�Ƨ��é>�eָ����ӳ�R�ι��u'�g][֤�y�Rj�ý���ݮZDB��,v?1j�ZF�x�׋WhA�7o��jN#�I�r4 �{���z�!�2O}�x��A��:�-L!�^���g̟'j�C�2O�c��q��^��������.�q�%��AC,nb�@�`�MpZ+ZͱQT(PLT�-�(ReC��D�3UՀig""b �0aI�a��N�C4��0�1MDID�Q%�)pș1�k�����<�#B�7	&��n.!Y�Sѯo�rV ۉ�[���2�F�ílņʅ�y1|�ZɝoM�.�k��    � �    ^a��^�0�j��,���,u�غ+��Y�o���׵���{���h�Y<�cY��v�9�&��4k�D<�Wm�;�5�"#��!��8�L@���p����w1�y9���X�+��:yg��%��On��n�+�CZ����s��h֓�)GT8�U�  ����aE8�i���+�5c��kx6�T�1��HX�k]fH�>�/�r���: �M���|=�(���$�b^2��Ԉ�J�)im���`q:$K��v��*e�Ւ�9�
�ۦe53Գ؃�����9$4��||{��Ħfߍ��Dܔ!�_��[��rs���rL��7'����k����Q	F�6��:uZfj6��-���$���~�g�ڒ�]ƠԚ�h�l7'����uɝ.'���%�Zx�E�)�J� �[KL��tv�(�y˝u�Q�:�!�=��������جx�H������������b�|�rd���I����3���ǰø~�~>֓�:Τ�9͌0�~����k������Ē�~~0{҂v�[7���ٛ��%!n5��f��r�U��	�yϳ��8Ng��Lw&��=�~?kCę�6�A>u��@����a�8��q�U�\�^�"א�&I������u�����I@���L��k���S+$���X8�%F�m�!�1/S2w'����<G#�M���A��9 ��{�}�]Ó��:����ffӕC_��![�Na�7é�0ӥi�NT�z���ߌ�9����VFM%��M`�|��I����ѭ�-�Z7�2d9v(���B$�`ui���T�^DaH[ɸr4�n%0=��3cԙI���o�3��>;�rd�Ct���ˋ��hx���zÐ�������Z�;g]���-�j3`�T��޴뢪k��^ӡ$�j���3�qy��k���;� kދ3��`��%v�Sx��׉4���߬	QM{lC�Q�q�q>�"�Ƕ�g�!�Rn����'߳�7I�����5�m`�/Z)�>p�"�Qe��*�I��tf�bo1>��Q��wq&eU����r�q~��?~�/0|��D<�R���y��'-�yy�ٚ,_�`�<�����]�Wbp�v[,�����:��zD�$������?v�7�����~�=��Ã��F�nx�u��O/����鹔��\�3ߌ�W�)3x�p�B�s�Yc!Y\#s]<f�0z���G�	���Y�8�����oO��~���Hd�g�ٯ�p�%/��`���w�c�R��x���|,��M�/�誄��*��:� ��^��M�&�z��B,�>�'��4!�u����p�!�d���bss)A��/��q��P�)I�,zyW�mp�Ȓ�-+�!m��^��t�Øx#��d�)�k�u�[\�P�.�n.�s�8k��Ǉ�EKil�mr�E�f�z�y����p����ܥ@я���X=JR�{�o�;���5���fǈk�<��u�ψ6��-%v�"wC8��3�)JN��Opx��nq�(hӧJ��#���OA�j}��㻄9���!�߾�i��Π�rr?}���b�I��T�[F�j�[]Q;!m�&�Ą�߫�� �WJRww�ix��r����NH4��s�< "%^�2QDN:2`��&̋����h\3�3.�y!�RGؚ@�Ԇ� *�F�ewR���)����wW+��@�������칸�␆b�u�`p�ON��]���J\~Ϻ3��0K���`����~��R����敒�"$� ���ϳ�[�߂���;A�=����%(��u������(}�>>���3�J�y����o{�xh�@��>6�ʂkοW�)���Edd��Ϩ}d��Im)\�Y����"ͼ��s.}�}���&:���ߍ}�+���[߫\)Bu�9�<���4<I�9)�Ȳ@�$��A�������=�r\������kv�mV̬���;N�R�q]l[m0��u��%�j�"�q�rC��^�Y�wwKڽ��v
I�l��%�h�Ѽ��g�4�������$�O2i'�~�~�R�`2K����Ilm��z�o�u��i��W܉ڥo[��%��7��w%X�e��D�*7C�b(ns�ɷ�
 ܞ��#�I.B���]�;�,�1d���lp�U �[J�B����r����u���T����9��Dƽ�f��? �\o>γ߫��{�BP�����9�ѵ�ŽD��.�OV��$��t���dn"��uO�~ߛמ��>�~*���#���~�z�^�g�c�o��n(�-%v�7�t�oiw�|뛙gu��չ�'8�g��m��������ZҊ�t���k0/ZѧZsl� f
�3�Lbn����:�� '.�k�t���t���+�/���{S8�Hk���I�����:ofO1>�7a�;�SNx~)����$���q=�b�Tٷ�@��O&�.&���(�Q�BH�L�-�?;��i��[�^�=��8r"�U%r�i]�Yj&�o��4�／F��1b�:���oӝ�&��^W�q[j!�rK!!j6�����=���������#�]��J�ȏ=����g�=I7};�i��x׼�v��#�nJ�:i��x���V�9߾N���S��y��Ώ�z"���c�F�֍�k6��p����������ߌ�\��$��IiUU��v��� �l��l���f�u']���`v�T�     � E�   ��w3�[X�B�kX<��D��al�FyqVsT��銮ٕe��������;�Ɲjܻ.ι�1��u�q�X:�IA��ͫX]��$��9!6��p$cu��=�k��Ҫ��j[n�3.���m۶����	�Q� �"�v 4�4� ���ݝ[\Α�����$uE�ęoK��j ��٬5�6Z�N]h"t�ۇo*�mS��pS�<�z�ѽkYfmn�8�	�y�d-]L�/.�\f�.!nўt�kr��B;���w�w=z\�� \�PH���9�m��3��o�tw������v!$�7�u��i��_ }҂�Ud���k��(�Rs ߺ{ȮB���4�,H]�P�$B���/e:���[�*o�;��;���]]�Z6ꬒ�[e �t��*���^��2��k�/|Ұ.��]]Zz��Z��{Ȧ�"#�z�'�h�ԳZ�aS��<o�����Z�-̷����6�p�QM���"!-C�/F�@bX�s�����nGbj��X޴�����z��y�1�|�K|���K\��{�p�UT�T%rWF���@�ŝ6V������Pĉr�7��t��;A�.�N�V�����rd���mL͕b��m��>~x�f󜗅<f���DD��Wz��6���k�"�VB�-���-���SJ\(R����{תn�{��&Sm��x�6�Y���Ms���\��ԉ����p�z�(?}��f��{����R"u��&Ш�a����,�9�4�|���׀��
�MU �[IJG#�b�7M��	B����'3M��;�Sm��p)��j�s���qt�����Ul�:���i*f��$����~Z���{��Rm���M�n�s+�s'���i��6������ʐp�t7vgfo!�i��΋��j.N���S�����KޖH���Z�8�*.�7�;:��C�u]6� y�ަo`'�D� y�=D�g�Z�l���P���鷦�đ k1;^����D��Ν��>j�jd���G%�J����{[�y/:��jU.$N(��X`�/�q3�����#[��zh�4��`�b��v�ͤ9
����TjJ2)���h-��,#4�a3��gxo4x��&`�6:�s1��@Hl�Mjx$i%����ӎ|7�q� �	�S<N�6r��t�t�
���D������<��;ٰ� �b�i��@�b)���)�-����'V�h��=�]�Żhrz�vn�F󪩦�	�$DZ����������>��;eRZ�A��k(KS�rHN�����m�����}�S�{�7;.�����5�f#������7�彬�m��U�p�tp�g�	;��H��R�rt�TJ�����e�x�r!*eV�%�����kB��H�'#R'`��Y���S����ހ��9ާ�v��"f�@���&�3:�~n@��b��g�>������]�� ��u q�t����as2w�?{�;޽Sn��d1{Μ���K*��%�YeN����'���&bR�������T���m�,�܇��S���$��:v���9-��Y%D�I�ONM���m� /y�ڻԲ!(�U�
!+K	���M���u�c�Rꕲ��Q�MN�L��(Z����t b�ΫWga(W�k��Q4 æM���5
�$c�����fd���Wa��&m�'@&�-��f�2�/Ƙ:�V�:e�G9��u��/�F��;��󇓶��^��1ӕl�m� �f'j�@u(Q	o���'[��L�9ӧg������z��޿�>�wM�>�0��id��+"w7��s���x�(S��R�Q5ӧ'{ �z�M� /�q=���9\�rTIY�����@jKw�����I�����{�D%.6�sP�I�����v�s�� ;<i��uH�9qiMN�=�][n�3!�w�ڻ �9�M �f�򞜛�d�x�N����GA��z`{ާ���p��@|8d݀fc�6��2��IH�v>�pS����9��D!AXPRN3P�Td�7�z޹¢sC�E@w�j&&R��&������5SX�y�^{�K��W�Um�r¹+̄�5d��6ќ�h���q��q�����t�V�K�       �m    Id�W��V�yى�>$���m����ڳ���z�zۭy8���l�W�����	V^%zՖ[dq�j�ݑ����Ohm�@�*��lY@�9<˞.K)�Y
����tö�.��ۅ�p!���Eβy4���Gt�gD�r\���C��en$16�77K�dvI��gft��(�]Q+�I����<�P�d�rV╿���1\�fg1$��1	�P��{:��/�����k5��\�n�8Hn�l�.������aqQ�udC\�[f��7)�ۋ2a�.�:�׷�o��MO<�vBYU���J�l��u�)='z��d������3��@�1;W`��-c��:�.B[-��%D�����������;z�z���ާ��������@���:UR����Qj,����T����7��;Wf�>��U�{�OKr���齀zg�u\�nJF��W+�	 �Ok{��'�߮��M �)������orP��(���>���޽�$��OJIڣ
���IKr'V����D�I1z��vy���T���y=+�)QQ�]�v�j�M�������v��������=��k��(��V��[f���;��X�ñge����k���.��4 rz�vn�<�޺����w��o`uMv�D� z�o��8G"r8�0�N�Y��s�wM��}�EǊf<B���HG	F#����{��͉�N����6���e��}�o�
!z�Us�Z&�s�~�� �9��y`���pu���~s��o`O1A�Y��l�r�YT�^[܁�u�6� w���v;!l��W[-D�������;/:����s��{<̄���{�um��d�R�Q�������ɾO���j�L�+���\�ɻ �Ǫm�1��cv��2y�Rh �1$��]��%�F�兤�HH���.�m���eڿ��ny�&�];^F]aRn�v���n�N 0��qO�ԳU�S���#�� ���m� �����~'�rO�׺�Ca�'"�}��� ��X�|�/�ô���m�I'�{����RX�ē�K)×I� ��xM�f:�� ����ROt������)cT���#�/T���K��;�f%�!%Dp�KK��j��(h
�	�JR�=&���io�^��z;:9N��!���o��ْ��>' ��ДE��DAF�c2!����|/��TӠ���3�ڻGV�k����mLO]��|)�W����]�f=v��=>ֹ��{W`e$�[��&�&�&�-%��ϓ�����r�
șqYC-���a��Bz�H�u�W`3]Nh ���u��fNE�~��ӯ_t�^�b'Zց�vK/��M���6��d�Ginz��1��:������Y�N��9�b$��`�pm��=}$����x{x�� +�<һs��(N��¦^N�(��d+���Kkuo`~bS��u9�bK�FZ�+�>�< �]���3rE��~-���'�]ĕ�U	Iim`�2����%��~���by��/9Ǿ�'�����w�Ԗ�!1��������*���5Zu9j�";7�#1�'^��d>3;����;�nh!7�CP�a0jr�V=M����`���F�v�HP�'�$��η�݀l�Ss@��<��=	D�Q۔���}}�_��7T�v�p8�f�efJ4�uj��c/W]s�c#�ٸ�Tz۴S=΋v�����#hW��,e$k���u{�{��m�M�9�*S�o|��]�M�k��ub��7�����}�}w��}��VbH�Z�*Շ9N�'��)'=�[���=9�75嶄�4׻��9qX������|�Uw�>�O@�||���\C̉cBx���i�Og;��$�3$��t��r{l���֟�B�����X܃l-�����u�� zs��� ,���Q��K�4�P�J�����ߑ= �\�jج�[
�e����_y�����nh��>��9�*FP\�#Z�g[ڻ ��f�n�SXDLt�f��x�6Jlr�n�@!���-H&��q��׻�)���y!�Ӱ�\�R��-M�39�dE�Xb؜�0}茶���������M��kZ����      $[@    ���\�F��乔�������JC7Fz�Ѯ�Vgt�=�'Y�\Af�@���FX�3tR6.u���.�9p�'	�d �UT�z%�����d��wlPr�yt<fv�8��\��F��t]�cf���y&:�6|�7��V;bu �u"�2��N	��[N��������ݢ�'.Һv�	����s���#����;@��"bx.�5�< y�p���f5�f��0QL�B�J��m��GU�l��F4��F
1bz�m����H�LF�2���Ъעm'���M��t����6�[���zr���ִ�]JeL�fy��v��6fP� y�8�N_�at�v�j*r��f�ԧP oy�ڻ ���Ƨ��!na��N���`��1��H�7#�&�Z�� ���v�>X��ls`� B́ЏɎ"�	��\�w�����R� �)'&�J�aJGY�{���N�c� �p���=���NjA5���"���ý���Ҭ�N-v�k-�Ҳ��AR�́d��xv�g�Ogꧭ����w W��9��3 ��U�̩ɓ�2�af�N�[��[�ا�3�୍T��wQxβ<��$]��{VBc}_;�ڒ��s��xѧ��$��÷�� �3��љC��1,���÷{ �]��B����JX܃�� y���K0a�3(sA���+���.����i9�yBQU���g㩊
�v������䩐�ᚻ"5	@����Nj���}����=	ˎ�IKimb&Q�d��zr�`ONj��{�XP�=�h5
�ۄۅ��� � s�z�O���XkN�c��&R�<ܐ���T� ~s��x�;�h�.y�˽�$��9��L�vڢ���r � d���F��;�I��\��ig�9����3�b�6 ��]Q�Y�XkMj&�[$����t�I��gl��2�4��g0�]������*z /�p�p��0��aFRG[%� ��Nsc�oY���b�]Μ�� �p�i: .����>x���:�T%��ur�g� ]���'�V��D\1E���M��,@�J�<$`����t���ƃ�<��g�N!L���$��*";�]4���bp�$�1$����Z��GqY�w��l#�`�>
�x�^�`t��.�ƹ�����z�.�>��@BQw���9��d���`}�'U�ۉ� ����g�6P
TGa5	��JW��͝���.q�O�,�[evQ�F�[���y� ��=�S�l� ��ᚻ �<ʔ�=30���[oKZ[nKq���8� תI-����m�
%��Gj��e�s3cPb]�l���p��ݯ8�`�Գf���ԡf��)�6h��Ī�����<�W��O@Y=�����pP~��
���imF�%l���$]��n�S̊�T�jS��)������s�Z��[ ߞ�s�9\��V�i�����[�̐>� }���eYJ�2g�L4�E�×{ ��ț��[�,@�d��� y��ɽ��s�y� 
��:�i(!JI%/��n�j�?Sݑ���uRF!wE�� �i�9;r�w������g��[�s y�5ћ��-���&���2�i��8HضV�cizMΣu��E��JZ��[�+���:\����]��Q��:���Ӣ�0��֬� �?\���#�R� �Vg������p� %��{Ȝ�8; 9l�Wz���S̹n�������:�������g䓓����ܒrؽ�v����RC�)z�1���m��������߰�v�2x����IdD�BN#@\�;��q�Q� \��ڶK+��F�T��Fo`��i�@RQy�:������n�p�u-�KM�m4Ѥ�j��~�y���9q�ݖ�e�,��@ �y�\�ܰ�eT�@��(��A��J{�]�%ZS2C������!8u���)11�!�TD
D�qP�}`ՠ*(���A)z^��+z�]1>c2�X�8Q�IL�[PPSd(�� ��.J�*�}��J�Юv� ���dҪ`J��<�@w�w�^-�0w�Mdb�n@ݢCR��.�6b���"DnH�Q��(؄��;� 7*�9dm	R�����&�f�0��&�	!-yYJId$AN�T(R�(R$)=���5G�j�'������7�_�;
@E`��p��Z-�q�w�ǄDG�CN���y�yc[��:���v�9/q��A��|�oN��!�A�h�L4�(uc
��$6?�N�΍�����5L�(�O��8���7埧�H����!L΋���A@@�aU�2�"p*d;^������o�8�GӖ<�[	۔�S?`r���تRݓ���j0��A�G���"(�����}5(XNq��̀������.x�cV�4�!d�V�R!2H�ɤ5������J����?o��!��@�6����wZ�V�p�S8�����}1ΘF舃\q��	g��~�
�6ю����*Hh�l����) T"EBBB�P� T$VEBdT$EBP�P�`T%�P�EBdT&EBP�P��P��P��P�!T$FUBP�P�!��H�JP��W�p���U%��Uh�j���)X�5�<Uu �*R�D�A�$tbS�&W�P��J}Q9@b@V�T��L�g�a`�4|7���b�#V��"��(��A�	�dP���]7:���{P�^�x9x@�}��[7�G�q&��H"0��b�W:�6���i���}��/�����w`�X��� Y��Ȓ����](2WX���2�֚ 7}(bV}���m�`ڑa;R��&�a"�|���	�����1�N�;��{0�`�0�DOHm>Q���x'�S��=T�'�p�آ���jj�ȁFBVx=<�=k��[�����XE��ڐ��X)��A@���"��[�|��l{�|�1 q���B�{:��2�ɋ �Vz�l�� _� ����!�ؔ��B�6Hg>��(_\Ȋ�K��L*8=�b$��&tf�C���Ӱ6�ʤ���QL2@�Yt\R�v��H-naD+��S�,���aĢ��	M�,���,Ь�Dm���w׬�ѥ��\䂈��n��(�k| �Y���X׳x� ��tu����}������>8=�S�T�C~�;n����Me�!��O'��y�1�X�aSy�(F��DA�cw�2}���W�D	��Z;�Q��q�5 B �����vi��< @��KE
ĠhO��*��=��xϑ�פ��wY���#ɐtn}[�pj�;��L	2�y��'���R�*I��E�0bi?qϡ�p���	��'u�&��v!���.5����.��*:������H1AD@ɼ�ǈu��i1��`2���@�i�30��K�L�C�y��c(�-��ќ0X;b����NT豈TM��3��/�6 ������C��DKr��; �GIrT;H���>�'�o�(�������;0���>r���ボe+��2��/��8�i�}	��rL��@Ɂ���yM�B���.�p�!q��8