BZh91AY&SYAj&z �߀Py���������`z�����@  w�΁�CA�I")�7��=G�OI�j=M��A�i�44)Hx���4@ 1 ц��eL��Chh��  h4jMD�#M ���  2h���54�4Ѧ�44i���  J&�'�i2=5��  �r*N�U���=�EJ�5�7�~��B�$ �g!��jN2�P���>�i@V�g�-��ײ��/�2$Zjd2�2��e��,���m.����iwE�ʼ���L&���(1{�,E���]DD��C	6�R� ��Fia�53:��ǖE
W��I$��
��TM�0M�r�M��r�����b�VȞj��Bm��@۽�1��4R3���*B�	k���Qz�`㎰�C�VU�&����l��5V�����vz�`|� �	����@��	�
eTm�%�L�����3:�@BA�V���Ps�^j�����b�ۮ�q뗍�K�fN�%0_ �̔�ڴ'9)[^�'2]�.��_��(��6�Z5�$�DH�]C.�͛6�Sa����5�O�4�lfn�U�)�@=. W9c�q�"�]@u3R�� �
V�}�׀�����|S���n�U�bW8v�x�`sN��j�� ��C��0&���W�(����XV������T$5Wh�1��$R㝛��ض�Ǹ��8L
��lH�P�`�.��ٟl��-�d-ӛ�e��lg،|�Uw�=f2oohx,���ɖUaSu�qp�Lck��Z����H���d��s"n�q[nE@��ъ0��UY/�.��j,�ݍͫ��� ��m���u�.m�ĕy�b�.i�Pe�`�l>b�ؑnڡa� ����	O%�ރ���������3�"O9�ق_�!����j�Uf��p�C���n``� �V�Gr��#��;�2�:���+�i~qNSr�]��@��UEE�UVF�v��~��iߗ ��(�� ��Y`ÞF9Ka���̚8*�B�����2���`�5P�Dq,�-��*[c0᚛	$Y
Rɛ!���%I�X��
CFp�&��H�D"D%xpHI`�ܲc�o� Z2$�Hw�}�kی-^�^u�HJ�,nQc�XaH����N�[*͜$�f�rtف�+���`���Ǌ[�ga���%ʆ!���B����f}��ސ����h@p��̇�p��}�Q6���yН'�@�#8Qc�	�<Z��B�o(op�����kۀ%�g��3���ؖ���
�uS��T�H	�,@�H�$D!0`��,��/�a��P+mI���t�8 5*$$�B!�f'^a�^o)膰�I�l�M�kr�p@o.�L���ll����Ci@�ĵ;N�=��:s���y�L�,.�������XH^4M9C욊�iȤ��w�����O^�0��˽"o���u��c��B�6�;�� g%!����q/�m*������@P�Ƌ���#��ۚ�\���WMZP�~��+|4�+�T<�Չ�z ��bk��;��9Xਞ��w̑�_ܘ��uޙ3�X�%�=4��O ��>3��u�M �9�ܑ���qTM��d����zv�qT�Jؑ�#�[J��*��J��8Q8�sݟfK�S��E�fׅ��:�TKsy��츔��N�v��F���x8W��YS@a�e��������tj��U=����H��seS4�W]��[)��a���P�J@�����"�(H �= 