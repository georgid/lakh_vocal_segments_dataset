BZh91AY&SY�J "du߀ryg����������`�? � �D4 %P �B�J���$�(�$���� 
 �)E 
�AB$E$D��(�)D��U�  *� �T.�   p���@�t)�;����b�@`�����Ѭ���7U���> 
��Uw}yU;�]UU�w���$Ъ����kA����Ԋ�� f�W�a�ݏ H�}����lԔϠ7%F�� 2������׷��[�@0^�����ӽ�n��R   5���{���}Vl4�=}��vu[�M�往wL�i���d��@<'������7n��r�^�����a��q  �4)�}:>�;&�u� =ޜ��tf^���wg�Y�c��ێ�
w�r���{��Zw} �'V���sw| ��D �h��Ϲ�}�1�N��Jzl�'���+l7��&�|4�����㛳����k}�=yc0�˻xx  �@    (  P 24��UI�i4ѡ�h   ��14L��RD�d�0�L�F 11�z�T�?RCM d  4��  Ob�JzjB�#A�i�@`�&F4�?B���Q0A�0M�M4d�L!HB$��i��&	��L�ɢmF#M4��z�}�X�a�������~�ч���P(�	�#��?O��
�'�?�*���EdB�������� 8v�g�?o�^~O�������BC����`|�g��������`�������s��-?}��a@|���"����9�z����2�����~^"  �f�N}'������>�gv|��=��.�s��n�vB '/��K��_��{����}����g?w����/��z�����U>�O!U:�T�"��U7"��Q�@7
��MªnSr���T� ��U5"��M��nESr���T܊��U7��M� �QSp���T�
��U7
��UMȪnSp*��T܊��U7
��UM���7��*��Tܢ��U7*��UMȪnSr��@
Sp ��%���!�}��8h��#_X��.��f��Y�e:��%8��U �Ë=A��m��S��^]�,Mj�[�#[����%:\1�A�rbI�&6�'F�8�'��h3H��%	�&���	BV!�t��	�MBP�	�%�$BQ�j}`��WIȪs`	������s1-4�y�v�:�1�ukw�Q�՚L7ݎ��Z #�����3;"��x8G=����8|i#G�@#��,W�cO�p���Xd�$3'5�;���J�	��)��	I��Ԙ��/^��2��a����:�AD5��ɬs�w~]T1����B���bњ�H�X���� ͐����<��J�V3���X3G�D
@PH;��-����c����"vj��n�îE��h�昋X��l�33g�s2tts÷��μ0-���.>j�:<�D�YfG�Pz��-o�s�c!�f&�o1�*H�
��XEb��R��6�փz�i�<�L<�u�r��)�q5	E��3��0�2��A����s�y�ힻ�F�1�{���k 4d�Ζ2v���2�ѳ�#5�'!ɩ"H�EfY�Z=w͆�'������f��MEIQ�:ͱ���N�sF�,��M1��dbړ��z��楆�
]�m�j1mS�wh*jk��G�yy&��,���Z�����w���T��fCr磨JS�J����2!2��%	ԧ�L��(J!)N�(J!(J��(JR��(L��!(OP��<���(u]&��޷�Ǻ46�(h/�Cߕ<�h����b����M׻Ϙ�|8z�ςmQ@�	`��fNC��掃zJud�'#%���'p��04;��X��k��PLx+�8�X�V6DoZ�Vl��Ys��l����9�&]�IrB��`+b�-���5���H�վt����f���f�t�"r1�����9Z�j:����ѳ"nk��kNjy�gLU�]�Fv�.V����͜w��z�:ٻ�ӻ��jӰ�q��2�5��Q�[�H��E�h�f�����ѷ����:�c3��3��m�F�=sA�\�z�7p���\2x��sF�m<ԇY87�p�u��M���W]�<y��f���wXӣY���乣Fa��n�S۹�A��0����4(;������o��4�h4�,qlR�x<STS	4/�ń+������PA�=�����W1ʈ�i��Z7țQ��u�����B#�DVqtkWV�um�0�8i58jw��V�rf�Pa6NC��fic-�$�ĵ�ѣ���N.BP��&N�S���h��#E�a�Q��N�	�ؔ����J��J�����jt�BRbdXHU!�w&�S�<�W'�Fh�I��[xn����"֍�ʯ[��������Ѣ���3N�͑hQ��K#N��<usf�h�F��!(2�����$��$��$�m�1���&d:�l�՚�Ƶb ���2-������,�UA1k[ֈ���g}��3["��˃FXi�Ô�a�^x���v��ݑI��J��4q�Оb���-- Ŷ�>y��N�g�x�HfXxp���z��v/$R�"�n�L(��	�0�t����7���u͜�[��東�|#A6Fǆ�Q[�@�,��C���/�>��t�c�^9ٷ���2����+�?r�Xxz¢����(��(���#~��:�����s\8���Ō���' �,�3�2�	�Ĝ���p���G�<����ֳ�g�`�u�XHP�F�4EKIi�C/c,C�Q�Q���0�e�d�k]ޚ�i��v�����5!�e.K��p2p��4�j���Jqp����s\��xuz��1���2�C���h�5o����e:A��V�fr��i��2���{=��p֋#���>�t)�m� {4��s7B����Ѫ���$;�Baдuh_�}F���"��{|4j%�X��z9^!yc�(��"b�/$F���us��zu��p���|<�I�e�j�9k��Hw����y���G��DyuC޹Nm���۱���������=NYbYPxk��ܯ
��^��@-Q�iX	� V�`h�(k��>w��+��^�h�L<�[ �u��1�N`bY8�X5e�Y	b`Yj�\oY���:�	�ģ#���Ԛ�,h�A�D�����;�|:*���z;9�I0�S�iȴ�ƀ��V�	
=ݞ�I������o����U�IQT�z2r�=z�cJ58df�h0v�$ ǆ�3>����_7gG�hK�(��J�_��ᇗկO+B��HrIn�I�ԇY.C����G��K����9Ldc&X�x��-uh���s��|�p�l��G)���4�#�wtz1�}aO]��h#}�4y����䍷a�j&��3n�͛�Sxe�����h�P^~t�h��P�4yPbǎ顺6]�%Da���q:�3[˧�37�%��28uN��\��\�,{��t]ΘѮa�gA���(�� ��� �写�E ü��@іî��@FFU�b���y�*70)`�J�f�B�A��(!j��.��Z���%��]o<�g7�Fh��Es�g�ni֭���R`kP�5��Z4a��j�O]�]o[�U�t:�e�����f�F��A��i��,�`j5�n浑������}=�}�Z�j*3F(���Z��5P^.�^g���{�����C�}ʷM���GA�wj��z7�T�����0с�����2t��[�1�vXN���V��2�f��@:4�
�����V>�״:�o�����@�@0,^,��f�zr0%Ú�9	����,d�r0��~y�%	JP�=L�<����{�<KF�2�L0����2ќ���h�'Xz �˝���> ) )�� ���X<��.(�4//<5w�����?�W�pDQ���7��$��Gx}���1��}�1X����k��,}�=��:��Mp�7��<�($:�4(,�mn�iUz�����)`�- )�a"�;ե ���03u{ ��F��;y�B��:HQB��ϝ��h ����(J��@��}y�[w8��E�6��Mw�rw=K�+�y��+D��&{&x��r�9�;;����,�P�d��>|������m�����C鯬}���ϼ�4*����~�p�H8�>_sꮁB����r�>�o�"-�Y����U*�>6�f����p �k (0��� )@A����� �8 p (0 s� )@CZ �J  d �R�$p �J  d��P�aJ`8 p (0-� �2$p�$X`�~H�X�k87E   
P ]�\�I&     A���䁶���藕��Ih jx]��m�HͲ&�Z浸 �`$[r��m�m��6�  ַ�� ��$  ��   � �lH   m��lm��� ۫n8 �� [vٲ� D��e�pQu��(���,�X0���r��k�o��%�8�m4��R���A�n��,�t��V4���s���\Zl[B�6�n�m�D� '@H0[=T9%��
�8�U� '@ �`�Mm�p	�����M��Y�ĕ�GV��i�d�U��-�k�-;is-� -�F�L�pd�b㶳c��m����n	mJ�ʠ($�mTYR
�M�   	               ��                                           -���g���������Ď$-�l(J����.Քi���e��6��6��  6�X��[\��H.��]���m�� m m� m�&�j���~ϑ|�[(���fl m$еҌ��[p�Y�t��ڲ���QUUi�rdP��|��|��/��6�����V�1�Vq��MX�%�ڧ�����r���T�ۥ��2۶����hMtU�;˃������P�ϒ[�E!ө�+Ղ�ne�$*��<�f�����lq��ŷr�[S�M��g���{��k��۫i4P��$��Ӥ�n���s`,4��ե�#��W�6]�MM[>a�ʲ��M\��YW��H4�n����	:N
��YQԑmy�N�	�f$��[A&�H e����^j����]thl����-���屍�_R��k��n`�W�eX6�� �N�Ӣ�fYz]Ӈa������7kh]��ڪ��W�uP\�+)�m�&�V $q��-��Yĵ�H��m;e����C)����gR�U�R��mX��%��|��Msu�[�򲓍�im���`8v�T��cl��B�;[�� -����I�l�:l]��<��)����[W*�Kj���H�^y�;�P[I4rv��  �iR�e����c���� ��	��f�sj�d�[I��S(��jڥl8U�������N�B��kM�I��m�:Ľ�x�'m5^��ݮ��@�j��^�k��6*�]g[�^�R�r��U�`$�ۻ �`p�k.�N�c[ ��rmd�3mmα\����|��1m�G�P�-4��H kE� q"Mm,�E�a�i���H��@�BU��V����Uj��Vޒ��v�X�۶�U��U�5�p�;XVVU�������)2���5��&�eK��  R��C�mq�ŵ%����t�*���r�*�\� �n���ͤ���rBM�6�Ŷt�h�n��6j�V��T����r�� $pBFĀ�K�ٻkhR�a�m�ږ��8mMGUZ��VZ�ڗb3��I�m��f�m�8���UUF�ۈ2ޭ���\�	~����mZ��&VV@�Q��W2�$ �/ �c ��U+���򟋰U��o 8�۷�  ���ڪU�˱���@���]���	��d��P �lUTۣZ1�-+�N��8ґɮ�ml�9z�:����K��gY�[A�`�Em��n؃�G3�9"j�� ���+�V�6�HŴh�*p�P WT�@R��UP
�e7I�6��e�IJh8��״�'HH�n�f��Å��_:g` 6S(=UU�m ��l۱N�UGS�N��5W]*�Gr�����p�`���<�{f�y�mO-���^v@���R�Q�u<ʀ��[m�'8��huX�l�]+��	sv�ͣ�	$-�$�Tی䅕ѻh�ӪS����
�q[�1)�j2��s��E����6��fVU�]T�Q�Z�[3N�lyi�m-�"@8�6C��`��-�k7m�&ݶ�2I�n�U�틲��@�m�qpH6�.K���[M�T� m v�t�m�m�$ 6�I w��ޅ���kk��FM�6����ӓM��� ���l��m,k��	�;k���[vl�Hm � u�v��    ڷcm�[�m؃  lr�krZm���0�V l8��m�m��v�N�j�p� �Cm��`m�  �k�l���m��۽z� ��6[Fεma��sl �UU���J�O�-��*�l����2@˝�5U*�����HĂ��lm� m�Xi �%	6��TIve[hUr�C��z�]���V�\j�%[v����F�;j�  [m�� 	6��Ŵ   � �mq��鬛l 7m��]6� pZkn��m���% �ں�%�� 5����!�z�$A���lM]�&�Ml�)�V�p �/3��
��˵һ4�WT#m�y��W(e�-��lhlְ  �a����ݶ A��$�6�  ��l���l k5��m�ۮl u�X�KmRA��yj�&�ymp��i{E����g�ۦ|�܄P=ۛck���0�3�F�g��[u�F�Q-Tp]1���� �CC[U �W]�]T��m��z����j�Z��iT�m�3�I�y�'B��z�O9���;������G���q�� � $��?7�W����[�H !�=�?E���>��?������?ǟ��~����* ��y��>W���_��������TR��@v��?H?��Ɋ�N �����J�N�h�P�zO���t �lS��[O�<NH(=��*l{W�(k	&IH�I��H)J�� 	 ���"��0Mzt�/����1��UzC�P{J/�����h8��H>�v��`���ht �N��6	 �	�8�T=	R�10H�v�(�,�t"�S�	⯩C�QBHpN�Nͦ+�}'"	⃋�x$��H!�/�]�� ��4���p��_Π�L���f���������:F���_gټ�x+��&���b䉘QX)@�&@	� � �%	BP�����*P �@U �4�.J�BR%!� d�Yį̬p �HjP�
L�3޾̹����'i}�z{�ƻ�.�l����g 2l -� d-�R��j�j�z�6�p囝�N՗��r��ܫ�V��EM�V�R�xը{r�1A��@\e�d�y�V17!&���T Z�$�E��]���YV��  �        .�uU[n����㮝��̃AP�b�фKx�|t�^Bu�I˷i<
��t�[�dM�'m	��6*����f9�G�+���
nrͫ����目2�&�`�z�m\bN3nn��$1��ҋn;��n҄9K���ֻt�����k�F�ح����g�D";uۏ+\Ʊi��T�<s^�.u�df	��SѺ�Z����X�Õ(+�&Wm[d��+�0�g����Q�K5p<�+�k��n�N-�8�ݡ{QaA�y�2N�61���F@,Y��!�j8��I.���8����pܮ쉺�@M�r��3�����Y�\͓��!��1��;�+n��qF�I:Y�X9"�Ȼa4�+K�Ņ���/ յg4[ I��`�Zuīt
3h�%,�TZ��\Ucd\f�+�b́T�Ut�P���/)Om�Z9c�.���:D������J1�R��9n��s���3z�{r�:��Y�1������v�tHp�zAP>��}��0 �B���]9�U2&���UO:x��Br@Eiq�D.usm� %�&�':�Lzv�ضݲ����Q�@8�.���hLs�g��75&7��F��ϩoij�u��ݚ�h:�hh�&v�x�4D�L���yNΚ�h����w���~?9��68��s��=������6�cz��ֿ��c<X�g��w���m�M�D�c��Ƶ�����N��rin��Qf����9�Y:c����!k�H�co�dَμw]x洒���@I,�Ι+[��w׍���>��=<e��*���m�sJ���.����"��֍�����#�W�����Up�<�0�լZ�Ɍ������wT���c���n�l͌ȼ����Wv�����|���kݸ�
b��b`�֏{h��]�~�����뎑GK�ݍ8�Z3�ܥ�t�/=� h�+�(��y׎g��t�{�+�H]�H�co�]dَ�O�^5�m%N��	(���|߁��c?g�`^U��iS���	*O���fF1Do���J�v.���3��a��T�Bt$��N5*8%Cuۋ�"��gk2���7�|���܍7�뮲l�{��w]x�M�T��f�t������^'u�1�H��w�Ͻ�B =�<�Zm[A^~{ӻ��O/Q� O!��e(�|���ʩV��;6���01j#���u׎��F���AT�7P�IN�U�=<��:.9�P2��F@HY��1�����s�J�yD"J�Ϲ����|�/���C�+-ػ��|�g1��~����Cۺa7v���c���g>���^K_UЫ�j�r�@�g�<^m���F��$��JI	R*T:5֚�)<"�:�Z�N� NT��~���)���B���n�ۓ`4�Tu��⸱�n�F�휜��C�]�ۮ��t�i�G.�����ҫt�@TC�YgFiz9Z�ն�Fa���6�{��\�u��t�B�ñj��za���w�|i
���;�26�dHF/[xζ�y�Z:c�ѵ��de8�:��w]u��]��r%�țx��&�w�x��ki'GY!f�t�������ԣB�v�) �Ww׌�o�]h鉓��"lQQ$-�֥g6�@g���:�yH��1RSD�qg�^7�:���Y�V�S�M�~ߟ�	R$�%��R��&���������-dԉ����A�Z<���|��RD�c���u��뮴t�{�ki6�ʋ8�z��Z�t�s�\к5�8���`sڞ7Wiv�H�@����nSQ9o�]hَ��s��n�S�*�X9|�泟|�����*�
ҫ������n�PÛ��({C�e������1��?g���F�Q�NA��﮴l�s׌�����v��>\���ݍ��m�Rud���r�m�RJ����$k�Lnm�=��{��g�bMH��w]xζ���֎��rmM22��7޺G9��gJ�:��WN��b	*O�ҹ1�� E5v�ki'GY!f�t�������N������v�6]_= �����c []ENuԅ�[kz���>�P�z��;aR�	P��y�:�ҫ���:n���r	�w�u�f;ܳ�|��/%υ�Wv�#�8��3�32<N��C�$#�3��w=u��9ȷ��u9ă �vm��� InɫL�h�� 5��ѭ\�>˻.�\���$�l���߻m���"{K���Щ����� �b����c>
%s��.{pM��ö�PVY�;W q��\��$������u���͝۔�t� ���	;.�����%���Nc|��g��Y��Ogt%��ҍ��q���  �y5���}�j�UUep��O�^;��օZ�J�c���w���1��?g�=��h:�w�~���c��{�<t�P�͡Ȇ�JD�7�&nlU�n��e�c=I<��m��1���=��zh8�QҒ%��倊`���|�g���C���R?}�絟��|�G６��ж��;���q֎��t���jF�6��u�Z6c���ߟ��������	�VJ�R�!q�fү$��ګ�j�U�Y�1���=��s�ZЫ]�R��c����_(	OJ��h:�w���{9��?��#B���1�E�-F�&H0�X>�f&���S�m`&�	$C2�!�E���.h0tGp�#	���H��0�xi���$cf�I!��1ݫ`9�V]�٦JL���@ԋ�oF�X�hl'Ya�Ĝ�0'�\�Fw�I�FX	�9�6f���Nsrq	���ĜĲ�Re����sFOȵ��=��;:ޏ. �O~$�v
��K��=��:�r���)@����!"B�>jئ�]:�B���߽�)N��JR�����ܐ�#�%Y!"BDȵ*��t*�1��4���iJV��;���:�~�j$$�`�$$HC�j��A�T�͊�ݚ;	"�n.������:l5v��n�R�B@����JS����4����>@7 iO3�Ҕ�'�Ǖ�k0ޢ��JG���ͩJP��ևp4�y�Ҕ��}�D���[�wt�:�BD����R��<��)I��z�R�g�yd��	�oUS�Z���Ȑ�ꖁ�)<��)N�߼ڔ$'�} �j¤��� \;�����w)JtuZ����k{���$D�0m  B>�d=�P��l{�tq��t�	��)�g7,��[.�k;��'&���R��=�ͩJP��ևr��� L�" ��P@�3�����l�k8�)C��Ƈr��~kJH��k�! )�%Y!"B@ȵU}���6��$$�6HH���ù#%;�~����z׽�)##�\���oĄ�H���D���;�6�C�z�R��֔�D��R��h+�|�	:��$$H��V}���R���ZR�����C�S�<N�b $�l������8�M��[�GKn�'e�f�"l� sX-���;o��\mb�����٧�h{������Ƶ��kvk=�8�sמ�1�1mqu����=N���]��iBv
�+@�(W3�F��7Z�a�a�BI8յ�V�nV�b�
���	��۞V��g6յwn�:��� w0m$mu�)JO]|hw)Ju���ԥ);��UNU7j�l"B@�&�R#PrO<��ܥ)�||f��(|��C�D������N�$�$$D���H�:�<ͩJP��ޗr��y�Ҕ��"��tXw�� �IVHIJ]���R��=�R���׽�	 W�p꺺NŷXHH��3��J�|׫JR���hw)Ju�S��(*�7�vt�t�9$MV�a�xm�[r��(�8�Uo�M�Sl"B@�&HH�ך�R�g�y�?擒�?|hw)Ju��[5�o,��)I��Ƈp_%=.fK	I�$H� bCr����R�����C�S�����s�����0ޣy��R����(]���R��>-)JR^������$�&����k�0/W Wj[�8�v'%%���m09�H�ڀ�p�\�:A�nNOɰ�;M�[6Q#k

!T�H7!CZ�r��(�ۀ���Z����9��v����$�p�Lk���q��Y �[��`�)�;��Uڀ���&�SoA�b��ߚ`w}�/y@�^�^|��%6�$��� �� �ۀ����ӺU"�K�ݍ��ճ^K���x�u���� Ht�������� u� 7i�z� �\O��I"i��_-��0.� Wjz��	����G%5����09��׼��n���wD�Ed���8�P^���_��LUcN�0=ͪ�i��jT��^� ���0.� {��!tU�-1��l��ӵK뇬T�����tf�B|�o��� ��r�v�ob�a&�So@��9� һP�n}���^\�ДӔ�������ڪ�G�� 9����\I."�(��^��\ ݦ�u���;�O��RH�k ߜ �
.�!A�v���dQ%5Y��7GVbq1�r[;lu�y`�� n�����l�4�rjuݶ�����4<,�8�ۓo�nY�ҧT0�iy����;X8e�6���7M�s�|s�rmĖYT�:,ի�5��i�6r���'HQ-�WZ=ߝ�=�j��r�ry:i$�!���=��㝵J�t��| ߓ�܀i{� ^�������G���w�4��8���n n�+B/v��dMSR�ր�P��تH�����9�ܨ���� 7����3�6�j v�.�D�ne6��Lsr�v���{7J��c�)6Zu!�hN������Iqv�[�����io� ^���`]�딸�� ��IuIW��C�V���K�i%�L{r�{�q��&���� ��r�v��8�w#���m�.ڀNn@4�� �[�F�:݄�8��}�����pV��ow���V�ӹ�m�Q�\�nF8`���>��_N��o�{�~ {��^_�=������&�#2�q��c�o���n@=�� _�.���Ne&��Lg���8�p���Ө��SNRK!��r�� .���Z��k�����^�J|ⴗ�  � '�K|�Ϥ�����D�M!FS"����؃����=��;�Ռ�2�r)"f@.������۲�r9*M6ހ��c��$��|p�U`5��������r��1Aw� ұ���5MJsZ������4�`o��Q
� �*�P!���ꤦ� �0ۈ������y� �� �� t>����	�������A9�yuЩ�1�a�ό=�e&�Ռg�{vne�|� ;R�Ji�# w�!A;��c��.$t����(��iX��܀k���I#B����K��rQ����w�6���$�M�ⱁꪬw}�@��ߜ(+���0/�������*%�G�0�;�C��gN�:Jw�3IT1��6l2��뮑m�0����7�r��b�����z�d�f;IR��aiR��p��z���j�[�:I��\)&�Xp�ցH�F&&A�\R�6ҧ�&��+Hd��:3"1�I��3��sAd�1���i�!�"h��6!�kC�g}�K@�ىa�&S�bdXA|kYs��㞄�}RIz�۷�6 
��p�� �cj[_`��6��CZ$ 6�Y��[M�W�sA�R� �*���ҕW�����;e����I�I��q�[k��9��F�6��K[u'p�r�ⴀ�Ɯ��e��ݶ�          �t˝����#���Ss��֎�v����@��e�䅳z��)�<eɼ��mG='.�y��=>�:���^�i,�n8=s�Z�f|��.�uѺ�:�9'u�Wc:hٹ�pdɐۭ���|��N4lu�&a�͙�<�-�Xpv���P')J0�$2�Y�2�`8��j�{͠*�݁��p\�ڜj�m�[)CG#�^�m�R�A�]�+έy�m/+U���%@�R܅��!�8��f8؍��ݰ�;��5-��=��\blORr������u�ua��6���3��( }�
:�V�{nܼ쏠ϗ�;Kj3W'Z��ç���"I�%��]w<��[J��r�:)�^U�"x�ҩd 횶��)4�"�mD/"�� �ܑ[�V�+n5�۞F�tF1G����3v�=���ֶ�&�8vx����]f8���h��p;�%��L���T
k��z��{fz6�ySyl^�KY�/C���_���w{Ч@*{U_Hs�z�}�˴�]  � ��6f����E���N^���8ؚ�ֲ}yg���u� ���t�k�icq�e\��t3��6��Bm���GC�l����u��ی��f�F�5��ji�e'gt�v�n1`�R��]��&)2�s N��n�nh��������}}k+���V;=��!(�������0d��3Y��#%e(0�������n�-�{�s�$�5)�hu��D���V0/W* ]��Rs	��̀_-�4�C6�����@
����P��o@qX�� �d �ۀn��W*T�4# _.@4q>�n�cf�>��B$M8�2*B�q��/'f�m���n\Б�Z��d �x�V0/7 ��S�b��6�$����	n� m�)\�@iB(��$n�Q4�fݤ�����"�/���oѷ	2�z��<�$(=�� ^��5����(�/� �� .��V0%�[�7MJ�Z����J�ޤ �C9Hr!��cQ�"9f��[�<;^q���U�8f�I�&�#2�u�4�0/>�cV4�﬷��9���_تT�k��?��o�k��ŷn�,IM�i.��׆��Hd�ҁ���D��|�ںϋU|z:�Hĵ��^*��U��X��O����4�f��Ec��07|�S�ԑ!6d�L�i��_� �� ֽ�@�t��`�&k�I��ƺ#�͢�:Թ��|���`up`����P�{q�EFJds����nPV03�+|q&ڒ-h� w}p��׆�� =㜡9�dfC����8�F����&+uU�}��� �î�R��So@qx`}U�1����>���o�m�}?Þ>�7
 ������u���d m��_uE��`��ːm���~�*���k��\���!#ֶ��Ռb�����H�c�����b�7|�S�ԑ!6d��ip`{^�۲��n�ni���1J��09����@�0#��oc�3Ȩ�@́�z@=X+�N���ix`_=��:���	����٤s!rn&θ�%�I� ��+$�ri���3�מ���F�M�U�Ӻ��[�#�Mwm[t[�;sqv�ŕ��nׅom�i㇫m�d���9�4(W+[�=�e��ˮ^B�-�ج�;*v�u���It!�E"���˶�Q�����{o��5�;����LV^�@��P��n*#2�p���R6�0=�H��O$|8�"�72�z�����*��c�PQ�}�� >������(�B2���\�� �H�y��X��U����Au����=�� w�p+��+ۺPm�n�q$F�a�r���s��yk.y����߽��jkZN'	Hl��������  <����DF��R�jMWT��W�ְ�}�	9����Jy�i%;�,V>��Xg8>�?�� F@��H6�B�_<c]��6�03~+|q&��ր矈�u�6�a�WأZ�� �����#r�f@=�8*�k�7r�v@5�_`7ARH����I2�h�#9N[\�Gc9o��L�����&�걁9� �[�UU _-�5ok���q!wr}��)V*��р{�~��0/ծ⊤i-hV0s����V+O�!�ၽz@5{�S��F����Ub�y�8�0'� ^���n��M��-X�1����Z��E��݃8�C����L���5�@��D�o8�*�ǐ���R�Wr�0`|pV0'l��D7MG�ۧ��UU�{� ��"�Hc�P��pR�wn����@.�0��BJM̤ހ�*�*�����W<�����U���)�5XǨ�V+>Ϝ�>���8�B2��@7�L�j�s�ӺUm��7����6Զ�H�I����բ�7� ��8s�3�xoz��wW�ƍUy��_�h�� ��c3�H��e8�$j�Y ��Ϫ���W���]||ouw�B�|��P�CF1XA�s�6���sM7�<�0&� ���v�N8*P#!��O��T�	� C;�����֍U{��[�C(	(	H+�?ߊ�d��%Z���y���=ګ~��uF.�R%�R�
x�� .�*����{������쮨8�M&4��IМ��ʾ�-���l Y6���u�t��z�۔�����0wT]���^۝���Z�V�c	Y��{u�Y��\��6e�Ʈ��þ|1����0��
rr�<r��1��f`��c@�D���fˠ� �ޫ/M��8i_\=b�ݤ�Y�_���"�H� C���kCNa'+ }�mp`O���o��"��s)7�-X���EfdV!+�z��y������^kr��F )P�I�pݳ���������0{��=ګ׳�̼����3���W�J���ewc�|�]V1�U��a�� �{)��H�ѐz�k�]���V5�2��"n�@�s����H�n�vv�^������ԋI��N)2�{��o���Rs��ݫi8��a*XSeހ8i"fb�ta�Y*�"�MkU� ���^��-CW�w���yh�Y�[�ۡI��9����q�/(�� �s�Na'ft�|b�����V0=��b�X���0�vE%&�Ro@yx`qc�pV0����+�CN��GN�ȜY���(�|�8�;�Y���qp`��V@�c�9\J:q���-X�c�S����h=�I��{�S#�m ��mpf���D��j�q�o�L
M:���E�&"�S��ӝm�$�����h!�fA�"*"	�"�%�a ��BRH	`�H`��%%�ffI����1�-���,�S��NC�F1��:M��AI$L��{�!ս	�a�	���"i�$d����4�rkf����&�H�=�PL�$�Y��1$��Ē{�<	͊�1����	�&:�Ց!4����w�|9w���P<O��(:_apUCڇ�B`�/�K�X��� ]�����8��m�?"�����yxa��� ��F�%Jd��w� �c���jI�X0��[YUZ,k+���*�b�&���e;���{�:Ռ]�@ʳ��+�J�Rk�����0��3 �\k��rj�8Ub����JQ̤ހ�cy�JՌ�n��wn7�����~�d�� ���c
��U����Xx�"�`v��58�Z��`��W{ǐ+����}X��O�����NAo=6ۍK^�6 �Q*B%�#Z�R��S#�CF@=�p�gШ�Ռ�ki���Ni���V �y �`{p��ap�T�f@�܀qpa�`.����`^��|��t(�z��`��
-X±E�� �9��0'#k }p�&�U�]����JI0`(P �������ٿQDV�n6e��@�j'�M��q���� �j�����7^л��L�{tr��e���5*Tbl��u��J�:֞<����mɛ�f\��L6���Pr�hݭ���8]�Y�K�O�w��>r#��El$`�v����fڬ�h�@�q�yu �V#%%T�U4����̤�@������P��r����7���&�M!^�1�|L�jǊ�`ރ�ƣ���v�9� �c]����du#I��!��0v�\!rX#n�ӧP;�x�>���Q �<�Q�h���]�T$�*"��B����;Nr�ˮ��]C�
uo��X,$�6Fs���2	�,���(����Ə}|a��V�N��ܿ8  �� �	 �%�iw��~�
�
�,,�/M�yJ�2���m�w��s����������f��fkG��0_��
R�0�0b���x��<L�c�&�M!e�G�� |$ `$wڏ�ƣ�s��VCgm��
,>��u�n5��GQ,��O3��o���}�͗`T���N������$gw��� ��[M�������1{�}�	 �{1��f{ա�X���}#9�̜����(o;t�N�������fmԫ���ա���9�)H�eH�'��܉��_W'2�Ʊ�+��ݷ�H��0�K'�3�仮���yT�����3�3'0o=�N]6պ�����d�f�>�K�:�.�U`dg���d�� D�N A)��ө�wUN��07y�������j�6���`�&k�>�]�q��sh�T�ڦFӑ��i�_m�3ǌݼ5��V��5b�O��w3&�&�Ȇ�v��;ò3ݬ͌L�䋸:vn��"O��w|�������o][J�2��j�3��wQ��R��qK�B���C��x!�[�,�u�4h��F �Q��XL��f˝)8�n�r�(1;%x���l�q�v�A�d�8��:z�h�&�h�98
�nX֮v�Nط@ Oj�h;Z�9L���-ez�L�v���H�>^�l�r�pW#���0�mc��|xE3l���>�������>v�" ��=>��R<6�9��ޡ��� @�ߥD����3�ߑ���<�C���KiLԪ┃ @�  �=�G��>D��Ţ��P�С�5�#�	"＋v���c�
"���T�It=�[�w]�ɉ��VG��A���J��&q���sO��*��A�@�@�=n=���J���o   � �+y�5��3"�޻z-�|�֟~���δ|�����
��7�Ϋ������L�%���<o\x�ӯ  @@ ����䢐T��Ƃ��361'��/���n�VثwUJء^4ݎ��f-���es�?~��@=����aUL̩�o��"�Q��!��m%�
i*�$�ަ`�z��9h��^��7�R�x$�{��  �D�B!����R�;�˥3�߽��ߚ%w'n��l]���3щ<�H��nͻ���	9���I�~�c'�ZM����(�*Y!s+9AR�Q���nL�g27Ds"o�u��3ҙy��|�8�5n��I�﹁'�љ����l;b�������L���ܕ3
�&aO�$�G/�a���M@���s��R���>�C�b���{~x���z7�gCHq���/#��Ge ]��ͪ��إmXI���s2k3щ���v����{Y��L�䋸7v�������;�`L��FdZ;��
��:1���F�5���%N'M[��b,�2�E�E���|`.A%_F�b@� hh����	�R\�\
h) :#5
L�K��a�C1W�NI0DicI�4N����dSP!��w�u�;����7o�$[��P��mJm[`8�8���[S�hְ�i6��/Y�<�v`.U��R�Z��-m�����I6ygH��F�6�B[]��v�f��"�����ӳF�r�hieݝ��            �:�g6�:uɑ.Z�ү6ek�؞�,,����x��$ �p<���lۓ�:�;���<������$(:ݡ�N݋!�61T	sGO��Z�N'l����L�b�KD���N�Q�g��y�t�p%����y�x\� ��;H�y�z��3�M7\��p��q��X)M��x-ݜۡ�.���6t�j�g'g��Nɚ�ey;�^�9����m��ɀ[�u�4*�.;ht��n��/i�a�������+n^��� �6�v��݃��N8���ͭ�˶��e5b��W���n���qʐ0쫋�l��[ˡ��Us��ػ��ɳ�<���Jndշh�J�T�tU+�*��H nL��K7�AeZ�ګjpZv�͇+��2*�T� �[m��^k�'e�G��ٺ:vɕ�zwdȧ&^���*���"u�aۤ٪����sێc&�p�p;�H�sS���SmͲN89�4�ӯ&���k����
��X���W`=
v>�WШ���ށ�;Ϗ<�����y��K��p���#�Iڊ)�p\4d�&� 5u��I�$�v�\��6�����3�ڑ=[<>�;����,�)Mpm�nܭ:�m=���ٻy ���t@�1M��l\7��:�����Ӧ!��U��F��.�c�:�S��$Bi	�Nu%8�W���9ͼwV񉑟}��ꓻUI�>g}�L��G�����)5�W�_��E���h��l-��4(D.<h���v��Cy���������v�=���bv��z�n�<ܰ�J���w4j
SP�"CY�,�i�
�Eqw׍�����ȴw;���Sftu� PN"�-�`OZ�)т�P@ut�H<K�y���gk>�D���uU�lg}� �Y��M��A��v�Vў�fz123�:�Rwj�:�'Α ���'�z1�b�^wGT�X����n�v�S�#�umrv�1"Α�"�э�fz2 I���hq!v���	z�����ƪ���*SH*AW����5�	Ix�|A M�=��f�b�U*���d�I���|h��̋F�UЫ�ʦ���g3&�&��߷���ۦ�m�i�gg>+gH��D��Q�ڮG����7��v�'y�n�b�U
�û�s���������wwM���'��s#Mg�^��Q�a�:l&�79�5� w�Kf����5b�$�)���fMfdc�H'};�պwj�Pf���gX,v��m�ԫ<Pd��2�O1Z�yA�<?�Fw��������w4��n�����{�1=�d�dZ6���;�tٛ��<��d�s"[��0��c;�̚��ĝ��]����3ݬ̌L��	� / ��WW@Z���n�f$��NfKs^�ݬ�X@�` 83&�h��j�d�vVsHY]`�Þ�ΟG!\m&]�wd���wjc�#]��c�j�tays��ӯ��эѨ�i�+vS$�Y��Z��S!D�2�V���D@&�����w��kv�y֮m�1�n-ɂwi �xr4E#䉰�ǻ׍玽�?�Kx��.rD52qJE�D�#�hɬ���,&�U��	��� ��3#Z(6��v ��٬̌L�䋫��ЧwUxd����L�D�����)&�ڥ�l�sD<	����*�u�Rre��{�\�.������.�LU�U`��O�hA �fo���$�1v.��2|�v�D���Ͼ���7v�J���;���̚�ؽ[A˱A�6ٛ;�̚̚Ͼ�ϲ���X�{n�r��j�����@�%���l�c=�̚����[�&.к���� $g�փ�G��J�T�������l�s�<Bp��Cq��3�h�]hJ�┃4=�#��� �o��F9�LU�U`���� �sO3=̐S��;l�uAL�ud���˥��DJ�(��r
(�**&q|��sl�F&F}��4v�j��?�H���֋�]��\ԉN�"k�$w5� F�C2k3}Z%�B�XI���s2k �����&��Iұj�S�:4�����^m�ա�3�ڥ"�Q�N6��vl3�C4�`����&�����L�-���*��R/`��wȻh�h�6"���wUX&�w��BV��lbguI���+�L��v�=��ޜ�m�M��2|�&	9~A�������o�B�L�P���W��g��ѥ����1L�]c  �!$i����wRt�#�׆��㶱�0kM'�㢝�ش�a9٨ͫ�9퓣��'�g�t�7hzCv��1�ES��m�m69U���m<�75��۸�{��ϖ ](����i�-P�PI���6�8���pV1}*��c��H̚���D��X�	<c���ȷ��hS�33j�J����Fw���S�V�]�Ӭ��;����H̋F�|i����1�ϐ���o����ݲ���ΰW<��u���	��+��������g�⊬c9�̚�	щ��9&.à���=Ў ��{�{�Nh6���3��L��}���*����m��	Z�#��n���ojT���S����s2k2sE�L#C����:���
��c֞��6!�U�`�A��<ʪ�f�x|$g{Y����7��û����;���ť#$$$Z,NT���#���'�.������dJ�� �\LHփEc3
pXqF%R#�X	�a����N���d�oz��-A*�5̴�X��Hs��3=kPIֱ]`L2��{޵�����J>҃�Px�A%�� ���}�.��q�  ���C�D��+����{6%�n���U����2k2swP䘻��>��]�3'123~S\��ɥ�`4��H닭�u����74��"�r2�=���}��L�܌}��m*���m�#���08���w8�)��!O�Q�Ġn�2y���RVnЧ�lg{Xkh�DR���o�݇wj�>e���OFfG����ݲ��U�NĖ��C�E�ܚو���'ώ��c�k6d���fdfMfg�]v�1n�`���d�d�= ��+��+�60�v��ho5��J�eMO�r���E���vf���ED.$���g}E�E�w�Hw!�
E"��=of�[�u�vz�UmT�!K�E�+��.#  ܺ*���=��w@�]��+[\p#͌���i��z��s��ݣ)KRoA�e�ոr=����zr���o`��'��4)��nV�sְ�]�M�r�@58듮+;�{߯{�|��S3���M*.�0���9�V6�A@��m����;�̜��1p{b�J���Ό�k3щ���s|�uwV���;�|��7�̋u*�A��tٝ���fMfg�]v꘻��c3��75�'����8�e&�4��B�QF�˛�7�<��;_;�3P���Y��F�ߔ�Q2����&O	� ��!��_q�Eؙq
�'��gF79���&�=����������&��z1�or�J�������x��y׳�����MD�IM��W��ݜ���j��ɯ&)*
�)���� /���S  A��"�fD��U�)myO��w�Gv����u�tŻ��63ݯG�"����1 ��+��+�'��k3##2m!�֚�bk�w��u棼�.�)��
H��z�;�kg��6�d{n��MPH��$�(�o���x����Mff�ʱWj�Ҫ�64��3&�$����VnЧ�:3���5����.}p������Ɇ�� ��ds`����� W֋�wbexʪ┏���b;�A{x�]��.29I��#�LD���%���:�1������z4s��v� "x�cޟ)�T\?��=���bdp�&�\�J��'����>�]�7�bbC��E�B���c	I����,+J�U�lg}�	5���I�	��]�P�Wv��[�x�9b�p�ZQ��k�ݐ  �k�[�i=ع�E˻zv�ۧ���c��ۮ���;SV��J���sr�Vf�4Y7
M5=#հ3�F�j2���k�We�z�T�V�@)5<ht�jN;U�zϵ���э�i��lX�]WuIа���I��)���w������}>�Wb۷o�3��&Fg�2-�U�UW�w5� � C��x��qU
P�S<�t}~E�E���3'�*�xgF{������ڶ'ή��%v�y+y���=�����%q�h˻uwt��۴���2|������g�KX�������p������̚����JŤ�	���s2k3щ��% �ݡW���3�s;����}>�Wb۷o�3��&Fg�j^����j�u��8�܎m��S��(dq�BY����M��n��3&�&�&�%�-�-�V	���fMfsS�ǽ>S*�R\-�9���f	 !
��^� �Y|z��@�41w1x�UDM��F��o5�Cؖ�U]+��3c�`I�b�Y���ذ���PQ�N-r��	f�.�d�'	f�b�m|����k2y�����*��x~��  �Fy"����q�)MP��*�w|�����ȷRo���tٝ��g��
��o۩u�i�wU�lg}��!'37n���'�@�m$�$j�(�$�G�cF.�ǄV�$��=��ɖ'�����UWWXd���123=��Ԥݵx�z����3=�Y����V-%}�:3��;5�����
f�
�3�;���c���"��������A�3��'z0ZTܦ
�1M!H��C.Z�h�6l�Z��p�Ű�8MY�	�YXa�߽���|}i�?O��M�n���82 R���� �چ@�lB���j�͛i.mp�f�3d�I���f�����@pHeZ��UIg�c�������+\�Ac�� +x��nƆmWT�{�$lsNZ4������඀           	]�M;v� b��Y�	mJ��c�@�5��]�X˽m4ѽ�]��[���v횋Z0��w`�5�8y���X���V{m�#N��/[�]A%��ɂ�D68rX�U��R%m5���bIl��,�R�c]=���y`�jV�DmHWm�'c1��Iwe��x���(l��d˶J�z:��ܙ^��N;N2���\5��p�o]X�v-�;����M���0�ڕ˗��G<�m�X�l�-��N�my��)��VA�y��k����'n�x[ass����.8k֭��H=>W=m�p,	����j_H#�ٸ8�xv�ۍ@��0��ݣ<���[�\��-�A�;2�ܭ!Rɤ"�Z�<sB�U��j䎝�B$3�0���E��S�(
{2��[�;n���km���c�ey;f����n��y��l+�T�T��A��枔����v�M�n
p�W��՗jc��׬r���mWc�	&�gA˿�ڊ���;Q{0X���}_�v>�D]�6�<bz�5����w!�Dm5P:ݭ�\�GjJ�/���T;n�>f,\�iyI�l$�#��+�>��e)��	��[P�G	+�V�s\�l�ܳ�4�ft�i�']�3��xK�5�$����_����������qXG���a��q�6�8diRJlr���$�;�<o\u����ّn��Wx�:?.�363�_� �?v�G�R�)T�ƍ������2qU;�l+�:3ݬ�F&F~�[ͫ�UWWXd��n�����3�)��%V��a[�#����vj݇�a�sv�Ű����6����3����fMfo�e]�b�W�lh G�  	�@M I�	�6�g��wщ��*��xgFw������H��������wy������O�Wx�>��gY��Y�����A���A;�m*Y��C1�qs��*%�b�b��`���d�f�'��uV���v�6123���m[����7���� ��aRE� ޾;�Ӷ��E��
UTOHx�!�C;�x�Cx���sR*b�@��mf#�h����}}緎��̊C��5ZCA,a������v��V����k3c#9"���M۫�'��@���6�qw��)UĒ;�C9�0 �h���[�94�
U3����>��H}�	 x��'��un�mU�ߣը͌d�gڧ84혞����Qu��M���7N2EI�����9�]�������}嵵�v��3����������e]Z��i+�'0�w1%y����#D�Ѣ���P̞���7tz�yG�]Xn�^߫���$�9#�J����{p{����7����գUF�wlM�9Kj����8�K�  �)��i;iѣI��M�a�؜j�D �����F���f�(.���m���L�r�'[�z�Ul��;@Cŭs�pf�\91��y˫g\$Ӗ�H�lZ5�{��^۪��u2�a.�uN�R��)��r�奘RR,ǯ���3��1%y���i�wU�I�sy����������SJ�B��������Cw��mw7t�'wU��07y�9�������t�X�1���F7$�/�T�\d39K�Og%�+�g"�����A@�7[g�~~~>��1�J`OF&�Х!Vl��:<�g�H�.c����6jZBA�@K$�_�^h?b<�Q�4�U������m㶦r�L�R��~c�k3щ���.��[��2|����Q�����mSt�wUWLS�W9�N�t`ۋ"]���[t�����Pu�tc����I��=]��]��]`�Qj�̚��c��m$�Ut�cFtc�X~'l�G�� ����O`��nuP��TD.	$��|5~A�\և���4*"*xw5e����|��_?_��t�T�w!I��5��Wn����'F�Z(%P��};��su0A0�[�y)�@NDe��<��qh�ݺ��1��ƃ����oѝ�16�3щ9�N��RO��mr3ь,�
��ӫy�������IM�1�3=�ة���B�]�SV��� 鍸�q����ղ�ꮪ��,X�Xѝ��g�j#7յ�Ť����16�3ь��%U
�i$�Όv�#=��5֮�7i��8�o�f�g�2.���
wt��:1���F=D{탾ul;�v����.�b5��%��:\�-�j �� �:� a��Nɞ�+���J�<��R�xʹ�[2�c�x۶2ƮzLv�\U\n��ݮV�xD۶@SF��^����/9u�c���g����m\�	m2�~��|��&N���7��u�a�`y}�g]�Rc�Z��N�������z㯶�b�n��QÍ�$�y���N�t��1�3���n��'n��>����az3�1��[A	iX�XџF7��H��Dg�[Q�$�ZI���'�#61��+�t�X�g��G=����%ە �@�%)�%D!J�C�7v�z�����H���ua�ux'TN	6 �$ ,.����H��'������������x���;��R�q@�S8'Fsy�ꋂ�9�TݧA<;#�`M�OF~���ή�I6�aՋ��g.�wL��@�����:�t�]��:0;y�5����մ h�Bfx���G��V��$�wr��T)�Q<�y���p��0$˜��;p3Q��k�C���		$Ah�;�:�+J#��N�0ޓD�@����טz�߬�t����`�8 ��}
u��آ��:� V���=�tuU
�iXvF/k�cs9"����۫��Q�bNg$bj[:��'v�1n۶�)ô�m��ڪ�
�L�`��;yWl7v4gю�g$�*#=�:��.����b�Df�$����mXvF/k�����mmWZwN��`��#��I�o�Kb����b�UcF{P`�@�z�[B��<ב5�*��AF	��N��<��a�NDD��Ӎ�ҕ Y��x���Z��C�.��Ȋ���`�������p}j��������1�}g�����]���XџF;�������6�WwU�H�o1r�3c[�P ���wU�Z���n��Ĭ�Bvn���<ۦ��ήl l66:N��5�]���c��n)�޸ƳH���ɶ�۳;�M]�t]������E���7S�y��F��b�C�� ��j�_�y}��۲�k��([2%��������{���﴾�~�7� �a�s8�R<�u�������LU�����ͣW9����}�;T�;�Wn�yIG��Rs>������.�e:#����bԔf��7v�ڴ�`�3��-IFz15-�)$ŕXgGY7ŋռ^�㵭Z A�iR��pQ��q�-V��v���������Tp\nɾ�z�  �G\f/MR	UJ�4HL �X �Fs��-��O8�b����`�Fw����.��ĞAw*l]���>�ǣ=%������jT���\n���z�z�Z���(�b�9ITi�TU�c]p�x�Vi��:�=�iX���Ό{y��ǔ�f��;�nڵ<���!pܗּI����������GW~a�@�E*��k:���<݌T ���$zu���m!�G\{����%Io�� 7��E�Ǫ��o���SlHe�(+$Z`�tuʴl6}�E�BHDѪQ=m�!�nY$�on�G�TػI<?��[�d�=#����´���)(�k��S#V�	KWUU�����fd`v�  Ԕoۮ[��wJ�V���c�J2kv�b��'n��t��ӎ}��\�́�9����iU�����1�FNc�3{��`��R���ݟ�H��mmq����n�e:2F=���ǔ�flM����U��f��򒌜ĞAw&ػI^]�z[��ޝk����8_Q%GRHE��gu�����5�b��m H�uZN�\WKgx�=��u�GE\n)�q���]��籺��Fے����n�]��v�0BpL��.�y7Z9��Sg�0ESq��;��(<��LZ�g��b������1sq��^&��7c�V�2i7��\	x�x�p:y,T}w�l���M�܌O-����)ђ1��܌b����-��]�b����qb�Q9��%�e$�����ŽFNbNf�\�ûj�yIG{�����J�{/m�\Yu�d�ڰ���nx��gv���|>|���|�Ԏ���rF-IG�؝4���U�H�0n p '�|��Dd�$��7B��5v�mp��{���_�Kg�H�^�_���$�nF&m-���U,h���Ļ�R՘�wco��dH����H�v��*ᜈgGArm�����l%%�����:���W�Z�mo��U��1{\�Ә�����0�ڼ���P$2�$���3�]��U5B8��u�F�Pd�֜�p�DύTԮ�^!͝���s���H��:`!GOF�h�=ZvԘ�H:j�RJ �&�B%�j��M����V�0ݪ����J=���������*��VS�$c���I ��4;�c�iҨ��(L�?4o��#vC �$@�tߐ��\�j*
g����o�{u{��绲F��R�$�qL$�D:u�����,��(2tk��a݇x5IG{X���-��݇Wt��'�o��������tҫmV���bmDd�bW$�u:i]`��U�A��=n��s�������py��=#7���k�$ 2x H<�RCb��l�df}NA�0j���%�1,!(�(��\����'�(p���PdA��Ӵ��B��aL��M$D��0�̒�$$��	�f98���I ��މ&"He��$a�`��@���"R	 �ႉ���"5I��i� �RkXd���@P4�!I8�aJA��L�I�3N�X%1K,㤴� CD��%X��E%�aD�A3C�����~�߳Z���v��A��  A��A�� ��`�� pm�:�i1uZL�UV�\���<���m����&م�Uz�8�J��i��,�9�7r��<�}���``�wЎ����8���nsU���           ;X�v�����$�+v.�lrƵ��vj�����(T�� ��s�k���c���i�^�]��p���n',g[�u&�6���=��mf�	�쫳�e�jf��B�r�Vzt�Xі�2����)' m3�ϙ�Skk�m���;��8咠�|o���gt;�=�-�8޹��uמWk��5'd3@èp[v�1Z끟1�\��waҬ;ecv�Y�[�9.Hy�T4����)H�y6�ZH��<��ح�)��8��Q����j�áF���<��f��t�v����<�I�n%ɶ,�����[�špJ�ʯ^�T=�]v=H͛<���	Mknz��t��S�
�<�(�2�*�k���5�R��RӜ
Kml��Z��2���ҭH�hx�Z�@`��h���mm��lɴ�{:A���Z����l��Ī�tFec��mK۪���J�Y��hu�
�3�t���a./\�%�=F������mw�����w���G���q��*� =���~~��}R�$)Eӳi1 2��ۨ�kH�[8� v�5���	.�<�k��HDG��Fx���J��8Д
]l�������)�q��ÞGԴ�q��X�hN�j扳��ek���iw�V�e�,�N,;b��W�ʖ@$�>����^�a�P:��OҺ�n�"H���;jt�۽���{���aF&�F�rض�U�X7���16�?Nc���	�N��F;k�������v�wl+���y�����k��ë�Xђ1��܌M���ނ�t�V���%G&�i�j�뇙���ZR6�I!�I%$�J�X��7�^����Q^�]_�z$∋8׼���ޡ���@�.}�A*����{-O fb���'��T��Uctd�{���F<�����-��*����3{�yIFN}}~~ߚ��c�X쾎�㗷9;f��1muqA�Gh�;�vu�*�,yoQ���܋GZ�l;m^��9��wQ��Ɂ�=��U5C����uߚ �%���;��Œ���O�Sb�+����<����{{�2�jb����2M�zK~C��|���|��;�(K�L=qll� 8�g�uK���ˢ�`ण��zF1d�MKb����ctd��w3r1�%��AƅU�X:Foy�)(��}�mm!;	�Hǖ�<�� `ReQ�3]
�0*L7"���ö���%�c�3�����_�q���(��M'k4��f���GR�������S�$c��R��͊�u�B��`�7�ǔ�d�>�Iw*�ut���D9�\�Rޡ�h���䠔T�)��4o��H����^��>5U��2F8o3r<f��:�)IRD�BH�L�S���-�t��a2=�֧Ś ,;v��[�*��W��o)q��ms;�yZg�8�n�۵k�6=F�s��V<�T�0��v�ɹj��on��ͭ��,7�<5�*,rb�]��K��R���w��Ņ�ǵAF*�WF<z���=��g�	�RR(4�o��G���I�ߐ���ɀ̪
g�����wq�F�cTP������163r3�[�����SgwP��kuD���8�ФUTO�E�g���[�9�bVT��IL��L�B� ,	%���q�	|xEjI]����U�>��o:BNLzF~�kz�N���a�`�@�@a�1=����;�+WH�C��2GF�C�L]ZRP&�)��h��=�Gw����)%N���F}�̜����=)��|����/P�/�qѮ�)��j1Ƴ��t�.�{���}��M�܌����ë�Tْ1��nF}#2p�����U��`vs@�@)�H ���b4�� �����'��y%é5v����}�̚Ǥg�=]��:�����3��}�u�y�����|�(�iQ��D�R��7��`��x��<�8�BUT	���װ�s�}h�u�JC�
��x;���Ϥg$c�%��N�u�}��9�c�0="���e݇xy�{�!��v �&��=��UAMW"[;#��3�>���NM�>��	ڪN������Ӕ�
����1T*B��5Q�����z���{|��Ԛ�J��3��rF=#?AսN�����=#9�Ǥflbyz��t*���ǻ�����3u�4*�u��gw����Y$�@؟z��]]UZ���&M��E�c�[7(��w�� �n�"�F뛚�I�{m�=��f�^��K�Oh�.�g�మ(�֕�����'+[�'����v���[�ڻgUP�:I� �G��P�X鉚J�G{�����V~g�lve]/O�z�v����n%�/�\lVѦlg���џHϤZ86����H�v!��v�0Dq��B�
��<GC����Ϥg��j�+��3���F-)�y.�5v��#>�f�c�3����t�:^&౱ť��\3����H��c�8\�������H��syz�k��]�m�H�$�O��ɬ��?�n��)U��#;�Ϧ�+uX���*�T�2a��瑦�����E��j˻xgс}�d���d�ϲ0��U��Y�u�C��&���f#;����Q���rW�Y��f�fNfz3�����J�N���3ќ�����]I��uXgѝ�1�@x)�(D�a� �c~�R[4�<FL���ȬL*���^/�  ڛ�A
�*XS��t�,#Y�!��aJ<9��)޷͏Ao-��l�;�)�i�3[���)R$�!��Fo���'�>�G}"p<��{I� �@�H 7�"�c�[Wu6���u�Fs����)Q��ԣ�b�l�v�>����G��M�6�B�^��ON�4�<òd��(!wUb��AՊV�W��Ϸ�����-�� ��+�=#�}�Ϥc�3����eݵxzF}�Ǥg�1�������6zF=�ϤcG��ĐȺq��Ɋ������g���F}#�w~}�������+x-,�L�l(7]�����;��ڛ:��#��$��-�g��Q4�����~g��zF}#�ԫ`�a�:l�{��HϤ`|7u�j�jت��3��}#>���-��Nº��3���c�2��w��ߟ]�>����5#��F����z�jc��� <�2Gl��I�]J���ûK����!`���:�%ɹ�a M�aJ��bzwj�N���6 �/2��bZC���,iZ�d���.rv������[@��uXح�qV�m�멨�_6��8��xcd�V-��5v��Fs��H����Ww];���6vF=���Ϥg�jO�]�����-z@Ϥcg�R�Wi]a�F}���Ǥg��]��:��W�t��s�x���ՍqGN*U#H�Lx��P+s����7FNٍm�E!5�)���}�������J��i	�mx���H��qs����7:&"U����{x� mm��suVj�]�!߿3��zFd�>R��ۻWx�����2s>������]ܭ��.�3�B�����&��#hT��T6��!����9Ǎ{�F~�]]LSWi]a�<{y��1���[��]]+��3}φ��$!,0�5��4@1*� �˹���xV��x����;���Ŷ���%!L3Jfx1�o:�v�.��^�dd��H�9)J8�ە��׋��(2[m�1Nº�'3���c�3r-�۫5v*�su0zж�o�l9�R����KfNc����}#2/�����S����G��u�0 �o���BTUDT������2y�H�OD�;L �t�mX�=J�mq�]�V8wQm�Wm:n��+��<C�X���'���x�$�=�̞g�3�n�A҂�uU��f���H̞c�kbA�v�a�F��[�:�=��eBQF���=#=�Ǥfde��Z�7v.ҵuwn�օ�l��b��M�����F&� 2^�\�Y�Py�Y^�����\58ܕ��;��9:��z�v����+��.�8]���9��l�<� n+cvSk�_j��̼�1��FDoG���M���Ki��뻽�v�6����G���5Y�Z%�$�u#iiS�TN��D�/v�[��S>��ι���V���g�3&�_M]YLSWi]a���2k�������P*x �ϛF��u�_�n����էx�'�{����H�xM�������@-��v;�2)�m2h�S�]l������y��Fd�>ж�$��N�͏�� w�B=���m��2�P�UAWn��hwu���q�����$��$Cz�2|��G���"�J�5U����1o|��~r}���7m)p�u�ϵ�82񱜢U��TXf�}���c�3&��	�t�]a��rc�32:S�xT�ui�:l͌{���h2��rFwۭ�uԭ:��#�7�����h��tUT�]V�3���[�ݼv��
U�iR��p�!A��lu�ń�z�f-Z��wa����163�F>R���t*��6���������!"е�:wuX'ў�3�Fd�>�ܛ��Ҫ�63��ɬq$1(�e�("EQ-�/"J@�͛m�E։�	�
��D�T��R �����|���s���M���,�N�x�6�Wo�u4ww
(�n��cV�	ъ��Ggb�m6�uA��Wb�Ӽtٓ�=���ϤG��̋��fbx3u2H rFO���n׈��/�S3*�Ep�h�1	�n�^�=���1E*
� �֏��u�*���R&j�	#��5�,��'㯍?���?X}��?�~	Ava%eUUT��"�h���� '�����;t��'����6o����vl�N�՞kjɡ��ZsY�E�6�R��)J�"WP��H�*(ĉ���H��� ����(��W%�$;Հ���D�/Ā��U�B��s��U�JAS�Ă������5�,Eܪ �!օ�MȮ�G�'F �y"/�"�(�b d���*��P:�`*�{�rU��E�;�Q����E2JUD�9"-*�BR �� �4)y����=�޳�ޓ�:�y�./0Zރ�G��� �R��B��R�"D�C�%|z��ϣ�<�}����/��0�G��Q��ؘ?�G��u�@_����nȒ?����I���>_�G��}�H���bʏ�����!�|����~�����|��4d@�>C�$:4|�ÿ�٣�~�Wf�{�=~��G��aϻ�6~{���������}�}8cҢ(	����t�'s�������~A�>�`~g�?��� >�w*"���L��~�g�>�������'�}���~a�~����p8?��+��?�����}J@�����������'�(��<�DP����[������?"4~���xw���v��ݚ������:��]}Y�����9L����Zuס�_�A�Z���Fz���>�s�:K��O����?Wߟw�����q����xn ��{ހ����ڊ ���>��GW#�[�р�?T������"Bd �%��$)
P)٘�j�%�
P"BA��@
d!$	B@�� $BT$%D !a	B �%d$BU��$	@��	 `!�%���$d!U	@D�$D	@�$DP�U !E	@��F �BP�Y	R@�!	a	 $�?v#�����J$*BBB�,!! H�)! �
����*) B���"�! ,�2I IAL�$!@JHAI B��$�(�����������HR I� D!����J*����(�(,� B��� �J2���I	� �A�K ��H������,�!�H00���J0��) ��$� ��� H�H�D�
P�D*$�(�zӽ0&t�ӝ}y�;܊b�_��C�@c��뢈S���������l�P@ON>�H4�Jҳd:��ä��>���~�����a�������w���__���������"��>���#���|�O�����~���}�������o���>x�?��"�p1>���c���N�K���?~~��g�O{����gf��u����?@���~)��	�L�����}F��~?�����?C��ߠ����O���ŏ�}�1Y��������9��?q����/�W����$���(	Ϙ��Dp1�����?���:ׇ�~����}�������I�����Fo�O�x��A�*"���y���XO��g�8Y?�3 �!��u��o���p�>g˰~�D�胤�}�2�`�GQF�}&��7��G_F`"�	��#�6��1�}���>�⇅��@|���*���5Y9P�����:�zd�<G9��Bo���O��_�������� ��P���w�u���������i?\���v~*��'��Ϡ��>��]�~����}k�& �M�����_�ߟ~���_�H�;�����|"���ˠ��?�f��jg�����
���A��4_�T~�Ο�=����I��%DP>�z~��? ��>��P����&	���'�=*"����*��ޏ��>����?y����}_�����w�dr�X|�����x���Ǵ	������z�� ��]�hD`Xk?�~_r~s�:���?G��_��~�%������/�ϟ�=�<'̷������_���DP�y���'�զ,2�Ӯ߷`|�v��w9f������7���g��c��{���	�2�~V���޾i�������٤�[��?��}�!������a�?0~R0��	�Y��F��M�~OF(~*��?�;����u����:>����?Wi�	Ѳ/�_��������1�t{��_��'ޟ������? ������*x�}�_z�Q����)��Q