BZh91AY&SY�d\�]k_�ryg����������`�  }ڀ  ��  h
 �A@: �
  ��ԅ�    
�T��(�)*UR�)EUP�����   (P,����_sv;����x�o}�/-�>��(�ضw� r�F��;��9�GF���  +�h��z�;�7 %@$��O���44��0�2��s�9қhK��8 GC�'���rh���������re�#�vr �
 �j�|u�����=���}ތ�kZ�� wF�Y< &C�7�=x/2ݸ��[�=���֍M���<}  �)@hw�ݼ��ۖM��}�F�N��:cۛ�j\4���	�ٴ��"{�Y=ۇv�������&|��  (���elz���@�M�}���a! {t�wWG�&�۶py�v��k����kU��9-�:�  �          CD1J�FF	��0�&L 0  �2���(�!��44	�2d�4d�S��RQ�F����bL!� bi�ت��� ���@�#F��?B���'� �  d@  ��$�� �F��O��3(��B6)���|�7��'��o��(�w�GȊ�cP�
>��"��A�PiT�(�� A,_�������4��h�_������/�����Y�=��V�A�����_�}~ǩ�����O_:�7���3P����%�@�*�  �%s(5?�;τ9RI%�ݯ���UT��"k�|�`�$Z=��뒽���~1p�{�2�8@Sߪ�t|)��������_Gˬ���_��}?��s���AA ���P@�!PPC  �DA� T�!�C ��DA�� 55552(d�!�C ��E�"2dDȠ!�PC"��E��2(�����}�e\����է���y��Vӓ���~�y�!K�!5�MHH�N�W[�ldݷiR�Ȁ�%C� }_S4� 'V'���4T
�L*(h�M�L����v���X/0��f��7E�lɗ��n@�J,1ԫ���(���K���NJ�������PYx��a�P�͚��D�Gln�$�@�\i��Ql��d�foZ6h��82�5�N^:�}��n-Y��J��B�H%�,�Y�N� ��;9:���HSp�L��k&/P)�9f�2앒kF�ͮd�`u6gF:��\�a�Is�Y���nF���E�;�7z�͒uw��G;�7$�v�4F����}�!�%�:�r	 ��$��N��K�UJB�(jPD�$��$"�Ph�(��5���)�4�A�DJ�iUoD��@�&BE�TD*��@��T*HI*�	���EWS��dSO}w5�6r���^��������*API�B�5y�oz:j�F�����c0�D�*�[�Qt\/a�Ä	p�FTh$�T��·˅M���`Y���*�QA�R�+[������*4��(h���Kmff������������V<���U9C�3\�0�v�����PI*R��f�s��8^�k�5a
�L*¬%�0��e�%�:�M��{��t�a!��.Y���d�*�0�Sf���%�F�c�]�C[Æ����k]���R�m��*!��.4P���w��}���.��*%_55(�\�Y��۔v�˘�)����Yt&_O����P���C� 2ԁ&kUHQ(�a���T2-K2�Lj���HB��x�;n��Q��M���ES�[�]�_�-�����*�q;.�y����j�p�A$�j�@):���hh��(
�D.�7��	�/��nރ�Q���0jE@!R��UB��:I�!u���uq#"�).��T'pI�A$�I�IKPI
M���s��$�,�\�{�GI���!0�eD9PNꝭA$4H�CaQt�q6r�4���ӄ G����e���p�2%%YS5�n%Ħ˙��l$8va.6��h�w� ���Ѿa��r�e� ^��l��h����37��t���tC�Ge͘�F��f:HT�Faѣ��^��Ѩ$�H��n	 �	 �)4�'!OAw�n	�M���B�^A$ ��$�I��Y��`�E�bzl*Jg��N��9
0ѳ\�oZ��/[x��{��j��S��	)-*A$Zj���G7ѻ[�H$�H$�HP�Ã��`vw��Aٳ',�:�}�sA��6��i�0 Tmj	�Q���
��$�H$�TA$E$A$뗛��ȅTF��	H_���/�$����y�Z�]$����I
,�35���.3F�ځM9�՜;2�z�h�,�6�-�2[f5!��7r�-�&�E�a��g2��µǆ�V��*�q��N܅Y�֋�G#c+���ٚ�$	UD�*	�E���m��<L�j	�'"��'"��6g5S�c٩�BJN��3}��7ٳ��th���**�	"�Pl*-5�HA$@,��� �.��V���Af���Y� ��sU�֞����p���QDi,�$�CP�B��$�H�\�T����7S@-�y�>�᫊���^|lmw�:�#��JK�P(j	"RTJ/&�T)�.l�n��A��0��n�N��d�D���6d(8ˁd
�C��%�+f8��Ѫ���1�I!v��S@zGE�S]^���(xtĚ@�)�#�%JJnCd�D�Ze�����2��D�]7tay
���Ł#r�HNSA��)JB�L��$�u�@��0�!j貂	*��n���I�����@q�I����W���;�Bи$RQl�E4ٹP�a�j�%�D�DY�/5k.%�9�х�:w!s�5���9ALj�´ T,���M3TBQ/4kz��n�O8��%R��	"4HHH��	%g+��K�fkN-No0�!*�ÃpI�z$&�3yM������;�.5t�*:�fB��SaT �I�W�u�}��׍��R�Laaܦ��M�̍XY�@茨P��QjR˧N�!!R��U���A����|�*!����n���3�P2uۛ�n��Cp�
�*\���8gS���F]��f�5VNH=h,��A;��!m�� �Pm�UQ�*�4I2%&�ӫ��cQj)�ø鑨$�dK0��é���p*�$�2/Xd�'8)4(�~ׄ��]�fh�9N�D�NҠ�*-5�ܜ�6p�z�Jm�fJ	dT�NF���D0�����r���j��.�R�3�듪ӷ;�ug]�9�%Kp�ST��E��ShU7#
��*S�����l�PHU.$.�Z!���i.6\e;�/4�Hy��!{n�/3�Qæ�AVI��(9(����Xo��Lh)�T��)�@a I��$�(�M���2q��M��+CM�Th��m����$�(/�E���D�BJ�H�%@*HFJ�Q�Q�@u�B$-2B��jA*	�	 �6B5
��ᠰ��J�@�9�k:F�pj���s'}�vo�K���;[�H$�H�p)�t�����j�Ί!�E�I�EK&8jv�p��v���)-�AP�uk*7t�U@�C*�B�����!#UIP��J�B�PQUPD�R�a�{ԫ�Ӹ�Էʢ�BK�*HF����6T���5D�٬��a��5t<$�=�I/�X�4��Թ�jM���cZ_}��y�/9�#~y{���/��6��$>o�?����?�u�gg���F��i����os��/+���?�}�P�}|�����6o�Nnݷ��o@ � ���mm$#��)�VE�E -� )	���i :@jgg;����ͤ�M�U�
��j
A�k��R�N1�,3 ),�i��$�I'JW�m�m�e��7Z��蒀�e�e�,�l��c!�z��l ���v�K��GD����Rq5T96	����m�E�����v�� k�-ɛ`ְp��� 4T�l�m��[&��f�m��   r�� $8[���`R��!;[[[WHMU3�m���l6��m$�p�` m� 6�8 p (�� ��         6؇0r��m.  �J �@
P`8 p (p82 R���t �J,
P`8 p (R���0 -hJ �Cѐ�pd�� �p\�2 R���� )@A��8�d �� ����� �p��� �� )@E� p��t �J !Ji0 $   އ�      ְ       �L      ' >�z        �  /Z��     )@    �p6���� �p �@0`8 �P )@A�����0 8`8 ΀ )@A��R��hH  6�_���������h0 8��+���>I���/�\mS`�I36�d��m(���9k]� %R�J�V�#�3)��+v�"<�~�W����g1n�R�m�]��A�'��I"N&�ͫf��jݶŵ<��pp���gvش����T�;Ua%�6eA15O5U�l�� �A��۝��uֳn�-��J�[%N��k���#��v��y��:m� ^�mp�PgR��.Z\1iV�@2^�^�խ�M��hh�m���k���d-ʁ�l�U]U@(�R���-��֭�m� �` �`[I�`�m� j�yZy��iv�@j��ծ�p�-��� m�M���5��&6ܮ��͵M��  �ٵ�ob�Z&�m��f� mo]"��lK&���0m�b�[��������[շm��JH 6�& ��8Ι4���i�Su.�œ�%��� $$m�6�Sn�j�{p 4�RB��kl$e�mHl ��hVj���^ap=[V�t���k�MP� �I3��b�  �F��6�m@۶  �&�����ǔ�\Nx�6�����
evU�/�nH�[R�Jd�����e�*�eZ��~?*���1�-THK��`��T8v����iLn\b�&�e�n@�++mҮ���+s�˴	9�55Ur�[VH-bս��.� �$ޚXͶ�m�Y( ��M)�����̶�K �0"ʖZV� �ηi8p �"�mp���{�z���`-�7���o}���zm�D9�Ydے[@�Gmm¶��(
�UX*�8%�'nŵF�	8   � �`6����j��j������Ke宫��� ��d��^ed�%�@4�Y�Ip�h-��
�J\�m<��/2�l  Γk���k��k����d�뵰-��,������� �6�k���������j]��K-m�۰d��$�`Hx [Zr�m��a#�� m�m��s� 4J4ـ p^��Z�ŵ�m٫`[\ -��y@��׶���	a֛n���g&Z5;-׬��e����{ 8��n����m� �zT�
�Ujڍ\ܻ-:�p j��[�Ͷ;n�*p��*��
Wf�U�mc��cm�6�	��q�ΧU�-��T��鶟����lm� ��lHM�*ҭTʮ���l�6�[@��q��Vݶ�Fӥ���m��ۭm���t^)���,FBez��n��
ڝ��v�n�nu����ną�Hɝ���k�ym�કj�Qkm�6�   :ڶ�� ��f��nӴT$1A =p�UC��*�ʫuuU@,�6 -���	m��m۰���K�nh^�!m��R�	 V�e8kiV����Q��%���`$8 �f�$ ����f�uUm�]�(y���k9��lr�@��v ��h|D�m��[m�@VԫOg���ԙ��	!� [@,��Y\��h�GA�@ �c��I v�/2�@�!���5[u[i1�      6�&����vZ(8` ��m/�V��   *�YP l  	i�c��Z�V�UU�'f�M�� ���m�@R�uUJ��Z�*�۵��l�m�8 m�j���xz��ڥZ�N��@� V�Ip N�n8)\ZV�+j�i [@ m�!"��h�fݰH*����)V�����X�t�m�m$۶� m����� 'F�m�`Q�W@�q�x���T�Wl ��՗��Ԓ��Ι��d�ٺ���Dm�����D���^��`;i�t��S� �t�٦���m�����acm�l@H[Am^�9,�@R�N�*��j�v� �l @   ���ہ:��kcm��k['`g���N�O;m��UPmN�8ͳ<���d   ��  m����m��6Ͷ  H	 m�     h��e�hհl�4��;ߎ^��Sqw���d�}���f������PA�c��}_^}?����� P:�={{������~���?1���5��o��<~�"����Ї���ߓ�����O�}Ꟙ<Aq�E�DKsJ��GbE�Q�}���F��6�a�KzB!�"2#!$`E�	 �!!@ �		��"�I!�Ѓ��@��J��D�
���c����#B$�R	DQ E	!]��S��J��P��aj�A
T)D�mG�,GT��N�,���J�@�:�؊�QbP�	h;E�S`��. �:���p T:N1@����N��%È�ڛ ҡ@(u�)`hQ)R��P�=�ҨR�`�v��j)hC�A�����@Hā!����~�ƀ��(��
�����j!"2"\ �H$�F�� H��
�
� �|�@* H�Ȭ�)" H*� ����� �2*��� "�"
H+""�"�I!$�"�"�� �+"� Ȳg���7���%Ĵ�w���vy�9���*�;`��.&�tv�E�j�n:y��]9:ݕN C�Bx�W�׏h��x��$��[P `�����p�h�G-���mXJ  �
P��[\ ����cm�N�@l �� �d��P`p���$� A�x����DڌF�� ^��L����mm�\��5�B횶N���=�θ^�k]��!ͫ�gLS:"���;��q��k�ٮ*����M�n58:���ں��c��r�%�۝�v�3�ܑ�cb�sK�R�f������z�[�P�l���n�]nq�va�h�ˤ��a<��m�J��:$��t�fu�d�49]c��䈜h�[r4g�F�nmZ���v
�D]��q�V��g Վ
�ֺ���q�G[&�M|�j����M�I������Zɕj��֛Jx�;=;2v���f�}e���^ۛ�2�+�]:vڒ�Q�n!Muٻ\�&�z�٪�� MR�\�mJ��m�]ۍl�4<����I�y@��W9L��a�6��NH��kj!�r.���h��yu��;T��j��k+u�bt�ZX�m�D��$:D��'��cq](v��4��n�*ʽT�=��S�Ψ�s�>q��b����F_��=V��̦us�{6qg���T�/1Eu@[@Hg�++��z$xa���쓌���>���\��Vlu�-u�z< C&:g�N�/RN����jY�V��v��nK��i)<�u�Iא�:�|;ν�w���p<l9^ݓ�.ǔ� q�ؚw;��J���'�W�Y����c�s�K�����9q{l�:�����uhZ8@L�s�z�������������}�y�7V�]�4=iy��2�\o�[���~zߑ�>SJH��Ak�����d��v�����$�cZ�<��q����/w�/4���++������:تdc"D�֖�s�����H���y��Z�F�6�(� ���]�|�-%��̰�9q����~z�*��]x�0�	D���H%F��9嶲�F&�-	�*Rl$�ݳ�y�\�bj=b 532��}�y�7V�]�4=��s.a����u¸�6I�ٺ�y\�
�M� du��Sc�EYy�+擰�%f��>޷������~�$�&�"hR;5��:72G����D�54��q�޷�������=_N�XoЃjb����
�f�lZK���a��^��Y�bPFtu�S�DGM��	��c>�����$�"9r�{�,D3-�9g޶y�3v�]���]a��)Dj�d�Z�k�����3�D�DS�	�9$N��-Nq�~�h_m��\��L�n.ٮ���˃SV�[�r!���n��|�.ݱW��0�s�������j�yv"�?$S{�R���^������z۶�	��Y$���]����'��	�eBj��;t�AJ��SȔ�s�ݴ���������:�73��]���-��=��9b�v9��sqP�g�6v��i�۶��z�G�φH�>��C��GZ���٧W�Ҵ3hw&K�ޓ��w7���^͹�'vog�P.�6K9�l0������k���.�B�uJP�N����H��܃9�ME��330��~�y�3v�]�<����:>�3޳Wl�m�U�B�L�n.ٮ���˃7� �Zp��1
Lf��^Ӯ1��n^H�1�T�SBM�4���-���y׫����k��'w\j�ywa�]�Ր:��"=��k��-v"�?$!��>�3޳Wl�m�IR�fXb��˶k�f�l�ິ.T����w������	r���i�Ɓ�ⷸ�FFlvӮ����B�������=~�l��3���nS���G�{�j���}�
*�M�^��Y�bTgF	ث/#*4���++du��a�ʳ�ϒ$�Za��o��;n٫�}W�B�S
d��Q�3����S��F���'I�&��"޻��=o�ug��i*\�Ħ!ˈ<�f��o��.���)CA:=�g��hr���Qv"��8��}�g��7lP!+�g���ܧ33������7�f���70�P�a�����8:��f�{s�؎a$I�I%Rmi_�5/�^瞯�[�mE��"J(��w������-%s!��n��;n٫��b.�B��PGb��`d���>$��ڲ�v�.ٮ���˃�U�[܉�����y!8Ul��#m�Ԁ@V�8��������RN4��M������],i�;-gaq\ծ۳ԝ�Y뗓g��#n�\Z���4�w�Jv�q{t����:6��	��;��}24<X{!7Er�������7�<��y]��������Oz�����Vi�CFȰ��}��o3̏!Vؚ��Pf\È�f�l��f홻`O��!�Nff�3޾!Wl߸�+�
@�p����Y��7�55mE��"J(��w��`�������Xy�i�.Q���)�5j��E):$z�|��-Oy�{���v"��B%LQ����{�f��.vbS�8<�f{�o����uh\.�"	���>���*��D��q={�u�Z������߆W�Ҋ��D�uȼ�ڡЭ9�GsK0�D2���faѻ�=�3v��إ|��C�]�<�7�f� %W1�N�l���:��ƀ�SF���aF���{B1")R�BIIB�tJ\�2��r��� �L�*�f�2+��$�*�@aR� 4%B��,B��6$
�� %�b��vХ%@���D� ���:�mIA
��$��ILe���Є�d-�41�$B�,�5�i���z�}�<�D�Zu�:@e!���A��= >�bj��g"�|�RE$N���"�)���$�+
�^]ޔ�I��X�RE']U�"2&���"�E�y��) �w]Ux]�۽V��qI�yV��H���H�מ^)"��yc�I��9W����i������g�p	�YuM��E�'�{����9�9�I���RE$:���j)"��ujH���z����
�K��)"���^)"�}wc�I�uV��H����H��~y*�̼��̽)"���c�I�uV��H����Ȑ�1�!"BDWE娆�9��r��$(��ʰdRD�]X�RE&���I�G���XDc@!c�8�n��E$S\�	R��ʕzRE$Ny�E$!s��-�P/��R����٧�43�kgl�e�qS�S	��J���.�����H��^)"�}wc�I���1j)"o׫�H���.I�+
�^]ޔ�I�~�r)"�uv��H��`�$$HU�䐐":�=��e��]��)�jH�����Ȥ��y��) �ז9��O
��YY,�+4��H��ʱȤ�Mu��)"��,r"�uv��H��!�N��\%�w�I�<�R@d=0<��E$S�wjH���^�r) 6BV����)U�������I*"`��z��p�E��i�Z[J�����^\��*Ȓ����b9�M�N{\p����p\-"#s��3Ӱk�6���hY�l��;u�v$�s���]m0`l�햓;.��0�8�u$m�G>��J�V��l���,�F�1N�ưl�>�nJv�������)�{ݢ���c�I�uV��H��դ��BD�Y�I	"�/-D7)��S�;�Ȥ�ʴ=�QI�wc�I�\�X��I�>�ՎE$S����W�e]]iI�<���H�+}V)"���Y��5:�MP&��є�.�l���RD|���RE$�ݎE$Ryʵ$RD�~X�RE5�+	<�¬���JH���^X�R@=!蝹$D��V�M@dS�s�b�) ��v�~خ�V�On��&������|P��9w�/��/��"�)<��dRD�X�RE<��Xؑj) �׫�H���;�+%�y.��H���c�8���EP%D(�(�IT(RU�qN�V"�=z�Ȥ�O\�S�*��7�P�S�aW$��)��X���;��H��ʵ$RD�Z�NUs��S��W�Űw:�w����
W�������Z{v�L���@�px���i�	$
Dc�4�N݇t���E1���c�&���
⾨D�̧ 3��7xĲ��ۡ]���S�j�T�s���L���P}��k`�p�;S%�@P*�����^N+$�5�Jl������}UT��&{%@:�� ڿ�{)p��������d�U�@^c�����v�Ha�$9Lp�3���^@]�U�¶��)�i-�����(�L����k2�Ӓ(�[q@�02�@���̣���[�� S�����%��@7���j�i���� 7޸.b��UOZ����>b_Rr�t+�}�us� gS/$/:���$�H���E&�N��k�9"
P�. �i��q7�2�q@�02�@�8�]k)��oa��10;}�y����洑�.��Pt�����|�K�ϔ Φ�����w`�r��v�RK�- ݩIs�3C��{�ߔ �S1%y �8 ��oϿ�����Z�en7b qr��B��U6�h(�Ҭ��z�]f���'VϬp�e�v_L�Wb��nl�=�B����[j;\=��](l���>_|x5l�v1�V0���`�1��WtZ����G`���!^��sŨ~���u��_�IDj�d��^:�^�ٶ	N�\iM���SPrEoj�ϓ(;}�������P���Ǩ�k`{� �����10%�1,��6�W`�p�yC�U����s� ���(JN�{�ߔ �S/$�y��k�c�7[�W@����@�p\� �2
�����&S��)4HS��'X��ɛg�w&���"�ܐ�� ��P���0J�e�*^�$�y��Ab,
cT�y` W�os�̬�N�U�O[�0�^��Ԓ2����Pi긃/$ �c�n뵕�jH��U�{�� /1�1sw�IuH�ml�H.{�`ms9I𯯥uW�N0�Fm�
�.��]�Y95�')S�¤'�b[��6�&��|�\�Qϗ숣�} >�t|�Bt8��.���T�wɁ�>��|�Z��5�[N8�J�K�����T�p\� �\9ؠ�8��ܐ�� ��P���0J�F:C� �c�}�V���`�2���Mk�Pq���V�rY�ⷻ	�F*Ŏˮ����Q�����?j s���� ^c�n�++���[ڰb`v� �8.b�n�i.��m���� /�p\� 9����Rr�t+��8W<�10�+E���:m�zj�Q�զ�����(\�g2@�p^u��߾�5c�Q܂vsq��uՈ���I����>'��~�o� ^c�b�(R���IƖ���|�b�(�L�%]#!݀w1�:�� 9�������֜��`b�(Φ^Hy�����SPrEoj�=���W�����)-��JA~q��>�P���4P0��X4�F����/Z��XJ�`v���N�VCS6V�@�$�!U���@�;��%-��I#(��Ch����*�0��8e�0�5�HH�@�Mj6p�p���� ͜D�o�	W��ȥh1"���b�v�(5���w�stJ�}.�s��r@��I#Z���i#P���Fm�vn��X�ݮU�+�R�	`B�iW�)��J���M��n@��l  ��h����(m��	���P-��8 p ��jM���!����m M�  7  � �[\ 8�7�{�zR�Ѣ�g�ph�tK���]d^�����i<�ܭ�>r���y�s���1s��	''T�����/-������,t$�=��6�.�l��٥�ڋ��|�YS;g�t�v�t���7���!��,�5�;0YG�j�m��,;W[@^�e6v��C��#��[��//���Z�j�� �����1 /SL��+�,����gr���6C��=#Z�mu5d#^V��yh� �mdL��B�j�b��.��y��n��Xb(U�ʀ�R	u�"�O;�D-�-mv0O%]UX+p.�u�+�-����6ݬ�<=�8�b����@�׉;5���:K#�6��R.�Հu���I��*Ӯzڶ�z�[��r���bZ�%C��֧2]m��^wn��i��4+�ހ�g�<���{��5"p��m�1q�����
���u�[	�J:C�H�-舉���m�p�T��U� �l�A�b���+�&�N�N
k��������A����:`�ڎ�k�g$�ز���,�ۥX
�4I�V����8�M]�n�]�l�]�l/y-�'F.Q9�v��n
n�s͐z��Z�k�\��^�6UKg8�L��m�:ܵ�]YRef�e܆Y+g��� ����#����$n�.�5�;bC�/e.�k�r��F����>�� ����P>K�&�Ϙ�Ԝ��
��|��������]��5������P�L�Hy� o�Xƽ����V�L�� ^c�b�PAÝ���-����� �x�10&�\N��/6��t.�uy$���.N��9R%%
��5v�� �(�L�H��V��0Q�\�2�V�*�Z�ԭ�+ؘ����V�T��W~��5$V��>L(�y ��+� ���]D��m���� /�pW� s]��NSm� �c�HJ��1039 ��zIn����������Iũ�k�L���a~m��Ȕ��;:I  � �w\���-Ʊ��u��`������p�b���K`fz@�\7W�ֻ� 	�D~! �{b�K����j<���j�
;���P��n�d`n�emP9"�Ń��`{� �8�<2�M(��TBR�n�q�K��:u۲�Ÿn�H9"��`����@�p���x�.�EQ�����޸q� 9����S���]�w1�;����kUX��0'>��H������n��@1�:�$�p�[͙K��wA탭j���7Ƽ�1��u6� �&��o`�8q� 7�W:k*7Mӄkt��t���3���㵗R80��A�q��3� ��x@b`^�:TLM�w@�r��� �&^H��V�� Q�]� 9���� /1�7u̬���[ڰ����ϓ����.|�Y�B�$Uml�H}�b�(�Ln�Wx�j(�BqGI�ڤ�;3`�[�U� i*�J���K/.�I�WUW%gqm��ۍ�Jaݻ=��3���v��j
8z;iG		��ݞ,I�h�e��M��`��0��t7���7����ۄ9l�A��cb"θ�!v��=��-��5���
���L�JQ�%)�M:��|�\��~UV�� ��H84|��F�����w�8�.�^Hy�x�Z�5�7[�V�L�d>ֵ�h��8�~P�p�b���Ka�w� /�p�1�+Z9����Ft����� �c��8�L�H�DaLa� J-��[��x2S6���\D�7T�����*�3��:�y5P�w\��MA����OQS P��o��$מY�O9}��"����B�$Uml��޸{UZ��?�� ~L	w��:�ӡ]�w�8x�@baZ2�@.�h�m�����x@<UR�9r ^c�{�:��+��6�؞�Q�zK-W=�)���|r|����Xb`v� ��+Tq� �9ؠ�8��ܓ�ҭU ��?��Ɂ{���UEM4��b`r�HsUZ�V��V�dL�$vs+j����%�J �z�$�p�[͙J�����s���PrD�e�}�`U]����Z�L =H�O)�	$
E3��Ŷgv�!����T&�T�慴H�6���Hަ[�6�X��e'R�t��bUkZ�H;o� �����䆨��p���&���Ǆ �S3� f&Ƹ�0}�U6��Fb`w��10����A���� s@k�ަI=T���GC�-��ސ�L�� f	�����7�,ks�e&�=�f����eт��{��7|>��݅b`r�H�OZ�3��=����Т�Ǆ�@wɁ�ݐk@ouWԚ��%{.�Ń��H�L-a ߹4cJEQ�ͅkU�!F�L������z�$@#^�����Ru)�I]�}�`so��`<�d�	ac�0��1)��$#$� H�H {�ǳ������f148�Y;r]p�CZm��!�ڑm��m*�@J�.x�z:h��سy,k���Լ]{X[�x�su�u���us�{];�������y�J_��7n��{����'me�"����j]<�u��ݹ�7m�3Z���l8�n�s�:.(m����ֵ_�*�PKj�c�HK`~y������� f&Ƹ�0}�U6��`�C�=� d�y��$����{j��ES�Tj�����Ӥ�F����L�U_[��b��{��QP�;�����Z��,�B�������$��irx�00�QF�O���Ο~VևIE�?8�Fg$ �L	W�����Z�Y�[�6���6z�Y:���rɛUQI,�͕u��2�Z��z_�� }��@e�-"�&�iH�:���y�y�ͽH��B�T�4�M@YAi,!����C�� $
I��䞫�VI:��=��X1A��UZA�s�Ru)�I]�}�`qo��UUZK�~��]X������j��D���X"�����I�w.I�ٔ� ���\�q�'e��qĖƦ�D�"	 �ۤ�݆��}R��_���-�BeHjQ$�!O���{;&m���ƨ��L.$��2�]�4������$RAlj`_>>�ECcW`|��Z�:�� Ń7��=���EQl����r�!4�!Ѕ����yB�6k�IV �j�\0�^	���*P͝)er�*��%�	IM�>Y���Gg�(f+e�3ȒGRF�#"�B�v��ڭƫ(�	�pP�& �m�4YK�2m��da䐇{��wK BB�v�Eh��G�'�'k`�6tD�����Igr� t ��T�1N�H |Wp �x�ڞ��̒M�W$��𫬙��\J�Ń�� 3h�x��&�iH�4ٰ3� z���@1`���*��&�!
!��&ҐJ����;Q\u���ܟ'o�5)�B݀f&�@1a��kZ��s� �pk��Lt�	l�~P����1:�~�/������m{�>_(�= >Ly��9�:t����@�
}.�'�L�sc�@P#3�(UV����0�y�T65v��j�θ,̐�k\��(:��N'*[M��3v��ovNk6Y)��U69[Z��iE���qtaG��@������MT�;Sn�Ń�j�� ��ϒ��P��+攊�M�=� w���Te� �`M�0�R�4�W`���}&�Ń
��|R��H+�_|��'@���w� ����� 3��Z׽ُ#l�¢qڧ��.Z��yڢ�������*�:eU�1Ţ󛓯v�sB�N�z��ݛ��L��::;\lR���ϝ�{��pn�l�M#[�=@�ӡ6���z�*s����cs�[�J�	�Ӯ��Å�m[�f�S����"����u� ���l��s��$a�~���ĳ������<�0;}��-� �Ƞ�5�3�!��k��`}�� �j`�aD.�V��&m8�Kv�����A���=���F�U�JA,d"�^��S$�weĆ�d��C�0C�32�U/!����A	�IQH�}��X�F�����3�7���9#u)�)�����g*��:�ߟ�f}�3��� Pݶ+�֖��!�
(�u� ��=�g-��oܤP�"�0a���W��Ի.䕡�����x}����'Tu�i?i��@" � ���l��1�G�q\%�ߦXb)��l�@> "H��v>G���z���n�����^m-�B�W���V˰&�\5�,�z6]@s1��<�g��sV�ά�pfX�������bz:�*�zB����xԞuݬ%�UP��1<�j���Nؘ�t P#w��6�Q��\Ɩ�!6Q�c�B��b5���Y�� ~�k�y΋Oq*�]�m',��F�p�dd�˶>w������3:�#H)"I�X�Q���츕M��{�`Nc�����)9伽�,1���g�bv5�1U�y���J(�  ��+�h�����H -ۣ�.`��%ĺ��@:�'�ln�3��W# �n"`5&%Bm�cM���Z�v[����!���i�#��{�fs j���y:�~e;b�O���͉�CRs�  �Oȃ�{��$HM�}��Oc��~c3άx�|�M��K*�En�s����kq�������:���d�\PҪ�߾����zvc��9��n���6�mH�IkKl� ��YesAl���e��Wv�]g?�����κz�PJ$�N��#���t!�;VT����1'/	�U�y�tz����r7Z��':��òm��*�j�ݦ4ҟ�� C<:^^m=[���l��q=�T�J�����Xa�.��Y�y���;�Ub�b�-���G��_��$�B�� �Wl[V�z(k����d�fAh]ݲ�� �75���3�ŒH5�Q���kI��x?~������M�/�)-G붶i�	o6��C��R���/h%��베�{����W�
�s�>_(�a�BX=9B8 @L�@Ҋ�:�,����~Y�H�x�~.%SG/�Ɓ�~���#�R��Xa�.��c5�19���c�Ū-���
(�u��y�1��g����gh�@lG�\S��jmϗ��H���{��~o���=OM���lj7�b���c��!���n*���A:����u���gxw�!�1-K��݇[�΁[I��B�%HDb�@�
�Z(
2�  sx@ ���;�MsZX"D��+������Sщ5Տ(�M��+v1A H���r7|��X��}�'��p��ջ۪7/k0`��U;� �>/�g瓯��籎���3I ")QCy��//l�6��ݶ{�1��s� ��@� D ��[lL,'GoX�G��ky�w�߇T�Y�+4{(�+J	" b!Sۻ���yg��,��ߵ��xxUљ�wZ�|�{"��J�"�H
DS�;�ۯk=�^�׷%M���˔�V�ha�;fwn�<No)�����.���?>u��&(jz1y�0+d����� B@��N�]��=Y��-�su�U]�p���W����QT�`w�R��������U�Gk��s$��H�F��^^z��R���?Ju�����[�g�A����	�.��V��R>�H0H	�����KFB$�B��D
H��F�T�]EU-�"F(�E㯽sl5u�m�D�A0�D9�Wme�	^������F��a����٘1gV᭖�=�̫�R�B����\�s�p6M�Mj�b�jU  pi�P8�6�p����� �@
P&��m�v؃��B  -����  7�` `� �-� d$8��8)�U5M�؝�\[�\tq�d�'u�X�t��������'ٲ��Ebݤe�lO��v֍��ѠVBjAO(=�,�����oa� 7f�Q����/>h�.* �N��)��y6��N����FK�iVv���2�G^��`�ON��h�gr޹�fN�'(4+z�|��ԧD��HM�N-n�k<�L�[��:�:t��)Z��<���l��\Ȭ�e5;`8)��Q���v]���;`c
l�K. �Pq���(�V���s���4��9��1m�gm'^)m�l[4�'d��ыq��0�!��=l�g�+��;ce���]���Wi�j�5 [S��s*ݱG) ;J�]�y�\��(�uk��{v�`���`�`�뇉�f��2�Y�L8�w ڵ�����^���iګ:6�۞͔yX�W-�!�����w��W��Ĵ�N�[;�
P*;B��R��2]d����*�֦�x׮(����ƴ��@mP()e����MD�M�7k��:H�5>y6��ӵG�V˙��m���4bج�땞v㗕s�s���pk�r��mv�hgŧm��;<��(����T��,����;E� �o7��Xl���@4*I�:��$��J:�#�f��uͯ#��?�$�
w���4\�%����}�1��s��ApI���|��Y������_ǿ�&(j�9��m��R|�}�LP��b��2`V,�YS��qq��Ě�d���wj�E]�-�m�=sm�7=�%%m�Jkx*�g�M��$�T5��$�Sщ���JO���h��KFQ �R��K
�c-P<)P;��tc�\k!Ӯe�ͼ|�}΅	�OF=�D�1h`�������bMu�?N*��[*�MP�5n���;�bka�ވ��baL�ܽ3�Ϯc��!:�s��h�vl&����a����u&�1CY���m�f�	>uݯ򆧣��h�b�w%i���櫨x�H�Ұ��U�� �������(�a���;�Q�-��1�H������O�Īj��7�Ԛ��g�J��?r�X�)�}n�P�泲�Y$��&���-(R�D�R�7u���NƠA��*��b�6�yR|���S#s����
�{�~e�j]}#��}�s:�(sp%̴� ���׬z�ޱ�I� l���;	�jZ�B�����b9�u����Ӥ!D�En(䋉��&��������{�����ɮLB�!9�O�﵉�y��3<�
Q�����H =�cv��������}MY�jlc{�k5p����mK�	� n�_���GkX��$y�lʓ�/W���hU� ��(tAhw�Y��K��y#���6���\�:*����M��� t���7)�7
iN�"�4�����`4As�ܴc���/m9�[] �/c]�e�i-��G�klV��s΀#0v-����Y�:���t�vMy�y�U�O���D쑌"���F0d@`�I �A��B
���F�$!�$�Ed�"�������^U�+i��vz�x��p�p��䚰ն]�dZ�oV^�����b~�� 	��1���%̴��� �}�rk5���vٶm��:���"dc3�Ia��*�
'1���������"����	`����Cs��]I�O}���5�q����3���Q�FҐ�����Z���������u&�1CWӮ+(6m����(�$�z@�4��ʎ����ȅ��0�/*O��\h
#k�a��]�l��5C]�X�]}����`Mwl��S�����Sы��MF[6�E�H�2�L��n�����bݶ�"Ѱ�l��$u��\P��rEs1�*2���1� �qh��7|̎rll8�QC��{��xH> �#1��������X�T��H+sX��ku� Z��^^{�6��[��Vo1qCSc�iA���f۱�g��|�w��66��jin�	2�F/W���{ОBbT���̌ZH$�I�[��n�T9�Bh[�e��F/����uF�Ʈh0pjڻ��	#��b�!B�zAUTUAa�b�F��]�O+duB�����M��$�aݰ�6�� �-�wn��K#2Q��<GI���d�zF<F�bN�����6���,D��6��$ v�7X��4.��VPl��$u�ήGSc{Ѥy�L$�ʪ����:���{	��jɼ�LgI�}�cv٭�9<���nfS��n�N[5�햻`�2B�j����6�V����S�ꍎ�k2$����f�`�'S���ms;=����<E�����}F�U
ί=��Ҽ���u�-U�Z�+;1N�wβ�n��Ϟ� ���s��vEQ�`��n���[������	�O�|}�[��Y#����[Wv��d�� B ۶ku��S[�!x�NdC���o�פbNuc<���Xh��HCdh�ν#��ۅ�0�bn�F3��#�:͎��%����f��[e�ٵ��OF����%M���`᷊��x$�����u�̑#��1ӣ�Ɓ
�$�@H^�{�c'0(Va?Byv�����Ĝ��C��C�.e�M1��D E�wl���W��"�Z��짂H��s��פ{�����r�=��:��d�n��f�B�L;_;���~'*�wi�t����[#9Ռ�*(�A�VW�u��$�^��U\:�p��n���:�o����v���d� ��@Ab�r������E4:V�F��/V�d�t�`F	(���#$U-��)��H�"�����V�,$,X�H�bV^!�VHL� �����\@�6Z"�lRS�
X0U�L.���	[1*�k5µ�S@(�,��cCN�G� ��E���@v�/`(s`y�[;]z�_���x̟:��S#�c�"G���L����;�Y�I�ɣ��,'0G�\S���ks�ᮓ3:ڶ��Z>{���׻��]
�H�`�0&������H�w'^����&�8����)���^�u@L��#��X.�<���g:�`�T��(S��eX�"�Q2�E,����o:����:��
�%�))4)$(Q��/k0`�쫝�L�Ǿo-e&n�F;�פu2:��\VPn�ʓ�B�w:�zF=�$y�L$ӣ��{^cI+��n����R�3�(Y� o��ݱ��y��P�,�K�u.��cߤ�u��f � ��������$�UԡXu2�dV�m�-����FҬ�R��I�U.��Kvt+���'��v�V�q�D���i74[�ۏHp�P��\:���n̯NP[������k�8������Ļu-��'@�ô٠�H�{�kZ�W� �ݡ�	$
DU#��ѹ�۱�Ѯ�
t<�__��{��յwe<|��ξ���1~���U�����vs�HĚ�8<�_(�A��T����I��#<�q���Í�H�v�􎀙z�+(7i���^�u2:�{>��#dݴ�$�v�X;U6�ٞ�v0&]pf�f!KsD4��1�י�f�$���yĳB��JSG{�u30�Em��g��N`���&������H�v��GW4ĵm]�O�:�s��פb�#A�&[���4E����7z��b�C��Cɛn���6��s�'S%F�r8�&�b��oY�z�u�g^�wu��o\Ym*T���w�{<�du��r�A�O�:��ܠ��[5�I��n݄������:�I��	�8��d�T����OG^��� �o�v�<����Y�Ǟ�>+w����O�=�uk���~>���;��߿m���'�KV�ݔ�N����Sс��H�G��Wm�#��u���dW!FFCP%4�@#oY�[ͳ��`t*� �P�$P7��Y���2.5����T����=���:�L����?qĊdX�,ݦ�Y젹���m[\��v�e��>�g��;Z�.����m��r�DJt%{u�
���7z��9Ĵx6�7Sc��bMu��И��[�4�}�:��W#���Z��짂H���S1��9�ě����BT�Ӂ�u�E��3�m� �ݥ]� g�<HZ:�*�X[�m�ѹwi�]�[t�C�j�J<;5�U�u]9�=��ghu>�ܤX9�FD�ۭ�1�j�˷h�شGg��uU>(�r�m�q�7W!�:��Bk�)4�����������;6�M��յv߫�:��^�����K��)el�������:���u6�T6}�ϻ�>.���y�u�bs��F����5��7X��u�������f�H����� �8.��d�n1�n��u�����4vL�4�)�,��b�V����M��#��%��.e�M3��d�Fx�$'3�u���2h;jڻ��	�u��Y�u������m]���=#��zF&�W�E/�VPh���:��c�H�ɭRK�6��]�'+m���tu=[�բ�J�x۷����M�H�o:�G^��k����O��w:�zF$կ�����Y]#��`�ЅP��h0@@")���~���X����n�Y[�:�sc�H��02.����c��zGY#�zj0�ٷgclC'�cMIc�	ڱLrQ$t���C�5JH�7Y�z�u��g��Mf8ǋq"a��c�	C�l���?o�W�E(�+(4R��{y��פc�n>d6Nbn�F;yפc���-��x�����v�	�u��Y#�H��G�g��S�ͥ��亹�۝�H�B��-\/���������:�OGY���n�YS��w1=���B`d]ݼot�gs�H�lu�A�A]�*�l����lu������mY���F	��^������S:���8�DK�(@�F J��$(@¨"�H�z���\�:���	X�̥� X@R�`�pJd! ʈ� ��.����Q) ���p$
��������n��BU(�hR @��Ȥ"�9[����T�`U��ݬ�@+����9g]:4�v��&�&��%v��hM�	UkJ��r�k{M˭��[p��`  �p (�mJ*�[H0I ���pm�m�\6����m  �z��  Ͱ �t� �m�9��(Ȱ�0v�����^6m�ݺ�:�.�l��OD�:�\�㳳;Z��A�ýl�@9��zy�hö�8���:�Fכd����S�D[<�D��ʫ�H�%��U�=shN͠GO2�ɭ�ĥ������:��c��ELc8(Sۃv�������8��<WY�mi�n��Ӫ�%��j_3�-U � �(���ӫM�!wE�rN�%�QS�֐^]�-�����9M�u;m��[�<�u�x�u���z-v�X+1��Q�|������b1��m��b�v���j�C	��%�S��Ed���hk���u����{�k��z�{])�X5넲�έ�M�4u��WmUmX��t�*��s�t`��5W��]��ɱ][ok�"6���]����c,=�;p�c)�6�\k�zwI����6�T�a7\`�vL�%@tuP��;	W�������Q@���R�5;�Y��U�����{ \�:*#R�Eme�U��2��������M��I�-y��vA�7Ä��v��x�$_V��sǞ��L�a�nh��6�<�5�v=j�a�/nӻ&�\��Oe�$���0�<C5��
��&�e˙��T&\P���^,�i��]8x�07j�����W��~��#Q����T����+�g���q�I!�K�z؀ݧ��~u��~�ζF6r����M�X8�v�H�H�0��#����O��w]o1�������1($�T��&s\ű�j�03�n[�8�d]ݼo#�b��zGSc���Z+3*Vh�\lH,�l�P�
P���X�4B	"i�c~���u��\��mu6����v�	�^y������׷��{��h֔�d6Nbl��w:�#�}�}��~t��Un�8�;f��х��*d�K/���׻�zG�l�\կ����v��G^�u��	������G^����D��@�i"���o^�Y�ߨ�4&f]C�,�23[��y�ŐMn�����Z
��W��~u��=#�1&�x>���-�v�\'Y��5�݅���DHôj^R򖟞�~~1���c�1�=�����}9��C��;��7Xގ���4JTP�}]�cH ���wXԗz����C۬�y�H�
�C, .�|( 3cbq��ݛ	7o+�c��HǤu3Ӆ��&Ք@`�d��vg���kd�br68�QR�$�n���e_z�:��/ބ�Ȼ�e^�?����Ǥ`\Ѫ�Wv��#�o?#�1s��n<[�R���{���c {vMs�������K~�����פaT� UZ U��%%�(��⦠�I[-N�j�qԲ6ŕ K��6��%"&��]���N����m�o�/�yx�Y���E�.}���j�d��N"���fp��٢���\<6vs�r�ڼ�V]�m�H;civka}k5^6���/w]���5	�m[�;b�/kQ�F.G��H�N���Sa�����^�>c�0=	>�7i��G^�c$`zG�Jޮ�[r��s.��^�=]�c=�j����`�����&�^���B`d]ݲ� ���^��H��t�B�E���4u=�=�5�v6cq�H�A����Rj��
n��꯽z�c�1sѰ��m]���;� �*�KT��$-+�B�0F��E��"'�_�Vkvz�Wp�y�qYA�V����>���1<5�/��ee|~���u�����i�����׷����{�Ct��vҴ�����U�6��V8�șM���l��n̈́�������blu�O�"���l�a�btu�^z�p�̹Y���,�Y1K1��%4-( @($ �UP(U"�@�P�#A���3��':;�D����w6Onح�7X�5���fڼ���{�����g�"fe���p/sv݊紸�Kl��4�l�v96>w���Aw�g1� �cz<�6m��Bb��ߞ��^�������i����}�׷�9�;����|ۻ;���1��H�x��A���O� ���I� ����ǫ�u����ʍ��D�ܧힻ>+{���-��:�
��"���xH�g:�I��5@�
��W�l`{��5�����Mu6�������bduy�LQX(4J�'�o12>#dbh��2�D��:Fg]{�Ě��苂��e'el�ig]ݏ�h�Rֵ"@!�/��pPR�˒L7fH��cnܜ���"������H��:r��J���ͭ����A&����R�Q N�����W����l��s99����I�qms6�E��N��"p�Z�J���-~��mg�]g]�uάvPmitbT�N��@7"n�w�2��u��:����|ۻ;���1��H���0��-]�k�0=���6�l�^zE�wv��c��zF$�M�Mwh��6:�oX�������e�M0��K��Bb�g��H=�p�X��śV�m���j�<����`zF&GW�D���Ph��O�4U
���c+�c�	 ��q6�m.�W ��.�׿F>���$�u��n��6:�sk�1��ϛw`�v�F;����L�nߡ��y]��N6�k�^�gx�9vu�����{[����'�w12>#dc=�b,�����#���1&�2h;h+�E^	�׷�P��A4Ӑ 1HKLbQBL.C%�Z����n�8��i/J @�it�)@��@��IeIEIt����`�	у 4."�� 2*���K�ߝ�V��HR����8 b!U��
���PLS �$N��=��wsa5�ڻO+��wk�12:��'���E,|���#�H�ȴ��msa�Wp���m��鍵]L$a���7�97k�w�F;9פbM`z}:�a7i��{��5׉���|ۻ;���ю�`d�L��	��Z�D�	>`gs#O�
�r�s��	�32�]��4�|�;�cw�wϟ[~o�(F��G�e��E��6l�e���l'f�Wh��6:��$�H�Ḯ�Sj�<��zUߘ�gkY��%��!@p�:����&GScFxkQ�"�F�X�c��M�I���;��v�	�״�k��J�3��mI`�)�q�B�)�\4P֛y�2jE���*�A+*g����]V	�n���"=�q�㭺#s����^��y����{�[���^M�:�Iݚ&M/6۬p���I�cGE��i�4r��hZi1<���5��S�׽��}��v���������+���-��4������s[�<i�6�B�2�y�ǽ�^�2:�'��j�x$��Fo12:��y�d]ݵo ���4ΌL���v�Wv��c��bMu��ld��Mu6��ʟF;���12:���$�aݽ��ύ�U+m/2Zͱ�vYLV�-Z�Ph�O��s#�� o����sp�8AM�׀x�$�8��5�c=�ZK=�m��.0M��y�&�2F>�y�n�I��T�1ݬ�����?@GWh��'��bf=g1�ݯ-`�QS�HJ�q���c73\ݶ�����2wj��1�Φ�$���l���)t3���H����n�[�lC��f���w�`�� (��x�s��%��!@pP�3r@��ZłB�k���[A�Jh���9�c3� �_ܥ�:K��hNHQ�JTTQ�'�
/="TɶjW���7��{�+u� ����^vۙ��}���`d�M���?@x�Wh���03y�60&�/=�B����6F;y����URX���wd��>��oJ��U��]�p@%���P$�)�U%�Q��:���mY0���j�v���F3y��z�Q�g�1E`��+����&�Sag�Z��46����Sc#>$��M�ݷ�/�|�f3���f�y�ndD9����Es��f:�c�T�,�l�H47
!؝n���Bʃm�QۥX

U\ڞé68�؞,n{S�y�G8�P�鎅�s��υkVLs�6��]i��'q�"n�[f�yk��u��z"ۧ(���+>�c���֟R�E�㻽Χ��v�
N��F��;<ζL�G"CQ�N6�{��%��:��c����H�.��ٷ�l�v󩱌��x>h+�F�	�u��d���zll6��Wi���o02F&�Y�D���A,#��}b�:������I5	�l���b��WNn͆�B��H�%���Ѵ�H�o?#c$`_ę�m����O��.���UeP���6/#��}<��n�$��*H���������h���0/y�H�Nb��Eڻ�6�H���Rs�uR�Ԩ�\oڃ����uSJ���ݍ��\gM�"�����vڻ��:��=#�����Sjͼ�>v}��ϣ��=�QXH���0/��:	���Vdu'1��d4f"������cGwd
ė��ܷC�~u��H�����7H�n�V�I�����$s��1s�<��]���m݄ۻʒ1���Ǥux	��Zd���`_s������$��32���c��@=��p����բ	s-K���}�1���GQ �/��[��՛yS�Ƿ�#�ק���)9��f���7cm.'R�ٗQ�.������=�>������u�-s!��S�F;y���H��I�֛	�O�[����Ɍfv:�����G/���C���	���B�&I��݃]�c;��q��WW^Ht�	��`Ⱦ�z�ʢ��
pP���Q	��B�"U��e�kCeD�D���H�Qa%1����
p � b�Ed�BF��B��� �A�� �`]� D� ����
 
��忆�>ݗ��I1b�vJ��O�?>(�	!��m��ݳ1٪��+�c<*α�v[v�"�K! v�.;�q2���PQH+� J�`8=\�J� p��G 2H� �J ���m�k\�^l �� �` dl
P6���p�$8��9�*�TQ�,�v\e���N�AW;�R���9�5�'t�
�{�֮�q����n��1�8'��fZ�
M���]�� ���5-]�1��ɔ�iOki���u��h�[���ѹM���;]FV.�%ۘ\��M�,�'pp���]m��<`�3r��;�b�m����␌����5hHN��U�Wl㭷]��H� �l��N��Vy�aX��� �<���`���-�ݶ:���.%�	Z:���ι�<�mC�tf�ΙL�zڶ�@���j��O\9;]�V�EZ��ڨ���� d��d'/EwA���-�f�Kл�-�ًm�f��H�	t����դ�����C^[��m���6��T�k!K�r�t].�]��2�X���]�����;-/��>u��[uYOFY�с�B0n*m��,b��y�l����v�@X�5ff]̄+2e��O��ؼ �B�@t��Q��O'R���r�:D�$h��2�sj�% -���! ��U�V
Yyu"Lj��N��gIzD�5m���e�:��+ŉ��5����؀�X,\h��$���*�M��3b�Y��V�.��n���}��wB�����S�w={��׽��f6�[�d����x�]��k�����~�"�]ݟ�x��s���a�U��`Mwl��>��{�'�5Y#=����yS�����_���+	�X4ȫ7��c���d4oU�1�Φ�NL�J���	�oEMٷ�y�V;(<�Zt���RJ�6!�������|��5~9�cv��-�a�2��� r����;�z�K4\��t<�`�|��Y��+�������l�v󩱌2*�L	�n�x'��o:�"����Q��v�aT%�s�.f�]�g�9n���6m4�l6��Wi�O�{�d�)�Ɵn�b��E�V3�f�c�����8�����5�X�|�t��P$�A(�G�oX�A������Cs�^:��c�EY#:�+a�v�я�r=py���Y�l �Xz��JR� .�]���;�3�<�ynN%1j�2K��Do16:����$]����l�v󩱳�EY�4����W��u��xȫ$b�a��ڳo*},��u�6#���Aګ�s}U���h������=#DM�}��x�msaWq)�[n�vk���]x'g�1�ܚ�'��?�s���d$�|�	�OH�w��VHćN�J�m�x8���C�U ���wY�	f�A�i&�/F���c9�����"�]ݜx�dc�Φ�<dT=gϫ�?�f�F8�K�mš�(�m�A�:ڑm�j�;J�PR�˞$9����ť�I9�9�dΩ�t�so;pj5������3Ӎ:!��f���vGI����"���V��zӠĪQ��`-��j�4P�.�zB����XB6pt
=!�4���S�w9n��ݿ}�=��I4-ݲ�Go:��X&E�T�}���o�T�K���q{�k1�f3<�B���@�dU��zGSc�ZN.D8SP��1�{��q��n�椶�[B�t=�΂	���݃[�mv!%�ahr�|�n�,�v�;�\Ɛl�۶���+a���O���HǤu�	�Ui�^2& � US 

�P���2GSc�}Eڻ������{�hѷ��񙡻�p"faD���>�:�d�I��i�Y���O���u�:�Ǭ��L��h%92)�Jm5&�v�f't�{J��.h%�>��y���2s4�_Z8q��gs�9����&s\�M�x6G\�ڭ�	"HED(�^yg�N:�+a��eIn󫑌��`'�9U�I��gA �����;�b�"��X������@gUΐ9+1ն�m�r�
�f*������Fw:���M����h+�E^��w:�\�I��i�Y�m�Iw�����u~�F(�$Z	eN��y����)����O��E���H�{�IΧ���۞��K�a�j�hq�c���a\vi��Ngr�|��}�:���F$<u�V�N�eIo�����u�	�Ui��T��������/=�Ii��[�^���:��OGY�NI4�I^	��w:���F<�
��r8�����K�r�S��5/;TQP�QۥX�*	�5�\�m8�ۈ:|���&�㛵k\ȫ��e�l�׫mF9�ɭ�٘�m�Fn�Հ�T�����y2����{[v�uͽrZ�58�ӻt�C������A�k7!mS��-��H �9�T�8H4&����&�����{�_щ����QXA4"(籑=��g3�@ �}�s�*G7]���s�߹��up�Q�̆�t������bC�_%l4��T�����c��z��;XRE�HJF�Dƕ3��͵�g ,5��J�Q0j��Zw�Yx��u������.��cD�"A ��9�g9���$�
ݤ��뻝OGW#v��o���h$��߭�ݩu��"FD��K*}^�#�9�����a$��4Jlݵ���vgvd����V��I��CG7^���u':�\:�e�!�+�뻝M��F$<u�V�MZʒ:��`��dmDD%$D�@�(��M
*� ��P$�-��p!(�D!
�Y��y�.�ˢbraz�8f�Fʽ���M@I
 ��$�.�H�,dh��c�)�Q$*D%T��H��B�! a|���EC��;S�4���@��U(�TS�3�3�ۭ>xuM��k*}^�#d�3w����[�^���u':�\ԉkq�ڴn�Нn���;�6u�\���I�n��I���x6G]��lur1'���|�o*H뷝\�d���H��!,��u{�d���=��\�h��ۿ<�]uo�ug$ �@�@zP	!�A �9f�\GZv�nTP�c>��M��F3>��<	�iZ�Y�,m7�ny]N���;7;eD�!���g��3��#���4\	I4Z����W��H�Nb��H;WwyozGY��Nu6:�l	4�I^��w:�\�I�`��i[ʒ:��W##�  VxE-��*�MYa�b�ٽ2�V�8t��eH��p[At�f��Z� g�:���㜭�`n"��Y��G2�th݃[!���u�N�ӷ8����u��C��t���6)9[�no,�"�Wn5x0��`kn�Y[�m�സ���Fe�0Ξ��:�lv�q:��2�ݛl[Hڵh��K�6:��2GRs�ZR�287^����R|�o>#!�26V�뻝M��F>��޵e�լ�#dn󬑉��2���d��::��'��9��D�a�-�mX�&݆��g�op;\����V��" 9����L�1�s��h I��<����K���G��_b� D@�AFBSU�	g�yn����$�0ZO��m�}#��:����<��Dl�+*tu{�OGRs���d4p�u��s�;���W�jD�N#x�ú)��>k=�]X�!��rN!��J��g��;�fs�'���,'me}�zA�:����+�9VrK��^[�uz�A�X$@��BA$����bk�� 9����L�1�s��q��+{��m��%�DM��]��z:��9r�i�EZj�'"k��WlI���k��@�m��v�o*}w��H��uy�LY
B���9�z$9�c{��Z��~����~���~u7�OGY���K�%hߝy��]����`�� D
�H�H � �ޕ ϷX�%�=1)�r�޳�y��c9��_���<�u<���\n��>�'q�s�:��G���ߝf�����羁 �]��u�1��Sc����I�&��h�x'Fo:���1����CQ2ft4�H[���٭�7ߝ^y�mXI�VT��7�����.E����r��^.��y�tU�Bڪ�DH�@m*�V
YyrI��\36j=s���m.�-�=��W6��KƉ��6��dVBi#�3JE6{H�']�M�0�/���Zu�l�U���7q�p��D�g�X��G���ws���'���\��`�w����<]����^J�`e�����{�M�����LE�!�e`�v���$d�	�j�	�YXg��o�d�OGY���U��/�I!m�<�����65��^���˩t�dc�Φ�S���ʡm+D����Bp��]u.	4�osO��c/Mn�W�6:��Sс�12s�d�6������ �.-��&��/Ͷ�&�YSc��|f�W���ZR�Ŵ�Sc�@$���/���Y�k5�� �d6,����|D�����:�3���i����ۆ��3lc6LjH��EIƷ��=r����'���D\��d��G^�bz:�����L̺�L�1�s�P�"��6:���w$���W�tu�Χ������ʻ�M�}w��H��u�X��v�4�Ɔ|�l�V�v^d)�t�{\H��p����f�����C�)k��p�u�1��Sc���#��V��Cf�	��{�"z:���zՖ�����}Χ� E�wd0� D	!"�4�H�K�H���ם=�u]ђS)'�::�s���c3��D-�h2��0F��S�@��[��j������2I���w�}z�Ǭ�fh^%�\˘t3���HB�l�u�� �[ͷj��0ۣ����gy�g1׳ѕN�l�L��v����u�GRɏҪP������̓;����_�>�����@��TD���I$�'�(���J?P �	�����mP�$By�L����FF=uѐH��+v�ՕE�#��T3�
@@.(! �� �R���
�H�"	?��*���n�EVE�(�"�����R��yj�r H�j�H)�C�BAQ
��2b����	+����S ��D�E�"
B","��-�P	dIBEU�4T"*\IEVDQ�AdUT	� ��QP�Q�YF�����=EE:���2 ��P���M@W"($� DS (��� ��+���[)O wuA��Ө��Dn��TW��{�_�P2"*H�����   �	$F��h8G�����w�����?�����	�G�G���oP�)�������_̟�3��~���"S���>�ϊw��!���%��s鳿��Y��������A���{�9@�>d�e�����>C��p�����?(O�l�u�tk����M\����|h������t����g������;��H��G���������'�R��	� (	�iB%�0��������|�'���w��+������?8�_O���ȋ��}��������У����A@I�C��W����	���#?����w>N�}?4���/�dZ�����I7�U�?�3z���E}�aM����@�k����c�Ӊ�_.�涓�==!��w������7�?5��L}���9 \je�_��v ��z��~�w��YB"� ��肠@Dp�%�@Q�#"H H�� H�Ȅ�F @�@�`�"��D!A�!� "�B �H��AHD�(AB�!R D�H�@@�PH!REFH��hJ@� D!"B	 "!"$ ��B 0*�B
1"�*,@� ���� (�"� �@ ��0
�@��"�  � 	"!"�"  �A�
$@�)b DD�A�"�b�D0B
	"
�
 A��@�� A�D 1 �	`�)b�$��
B*�� �1F(�b�1�B�@�1Pb�PH# !�`�X!�1H#�R ��0D�H#H�H�!  �B�X��0F ����"�� ��0`�*) *��"��`
B
$"� �*� � ���*�x��	\[����s(�G����y������6b]~D?���{�'̔ "v��Ж��U�9Ѵ���>�y�}M���J>c���@Q�^��o��Pd����������D�M���!�@����|?�b}U�����>;���A���b�(	������{;ikF{�������̠��n2��u�<����;��>��z��m�����x���ߺߓ��A���},�����������FW���K�>j�|���W������m���D��}�쌊-!_8}_]7ڲǳw���w���g��Գ��#���\!Y�'ϔ ��@��A@O�:���H�O����4~�?�@}�C�:dz~��8-0�{p�(���� m>�4��xܑ����u�lߺ�T������0�G9MW�����:'?�����49RH��:\ J�I _�
v�v�bx:�����Ζ���q�����`tZ�����((	M�M�~q��?Q_i��{ �O���
8}� �'�|������o���~?��G�������������㿏�7��
�q���}���H��������+)���>d��>��y��� ~���0"������u�����C���?� A@J�~Yo�{��>W�������0��>������A@J�`m��Y�~���~���h=����[?7a��#S�|C��C�>^��"A�x�¾���u�ވ`�G��x�!A(��'���|ԛ��<�������~@�ZC��>���/ہ���:'���OUg���ߐ�����Te���r�Q	Am��������J����}0�~G��=�r��G�^�=y>�B@S�!;�'ǻ�tt���{���~���C�??��ϖ����# D@O��>��0�D�ge(}����-s��_�����>R}������f���[�_��q�wK�0�?�M��o��'ҟy��k*�$>�����)S��͹������"�(Hl�.~ 